���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �_sklearn_version��0.24.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hNhG        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h-�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��h6�f8�����R�(Kh:NNNJ����J����K t�b�C              �?�t�bh>h*�scalar���h9C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK�
node_count�M�nodes�h,h/K ��h1��R�(KM��h6�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hkh6�i8�����R�(Kh:NNNJ����J����K t�bK ��hlhvK��hmhvK��hnhJK��hohJK ��hphvK(��hqhJK0��uK8KKt�b�Bx=                              �?�'�V3��?�           c�@                           @�������?�            �v@������������������������       �        �            @k@                           �?����>�?_            �b@������������������������       �                     .@                           @|�-蝉�?W            �`@       
                    @ףp=
�?-            �Q@       	                    �?8����?             7@������������������������       �                     0@������������������������       �                     @������������������������       �                    �G@                           @����X�?*            �O@                           �?l��\��?             A@                           @���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                     7@                           �?l��[B��?             =@                           %@�<ݚ�?             2@                           !@@�0�!��?             1@������������������������       �                     ,@������������������������       �                     @������������������������       �                     �?������������������������       �                     &@       \                    @�������?           ��@       E                    @ �J���?W           ��@                           �?�lb�d�?�           ��@                           @0d4�[%�?�            �q@������������������������       �        y            �h@������������������������       �        7            �U@       <                    @<ߎ����?M           ,�@        !                    �?��=<�?            P�@������������������������       �        �           (�@"       -                     @�"jd�?f            �d@#       ,                     @�q�q�?7            �U@$       %                    �?�{r٣��?*            �P@������������������������       �                     >@&       +                    @tk~X��?             B@'       (                    @<���D�?            �@@������������������������       �                     <@)       *                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     5@.       1                    �?v��:ө�?/            �S@/       0                     @"pc�
�?             6@������������������������       �                     @������������������������       �        
             2@2       7                    �?Dc}h��?"             L@3       6                    @8�Z$���?            �C@4       5                    @�+e�X�?             9@������������������������       �                     @������������������������       �        	             3@������������������������       �        	             ,@8       9                    @ҳ�wY;�?             1@������������������������       �                     @:       ;                    @8�Z$���?
             *@������������������������       �        	             &@������������������������       �                      @=       >                    �?���#nŴ?-           �@������������������������       �                   Њ@?       D                     @ ���J��?            �C@@       C                    �?ףp=
�?             $@A       B                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     =@F       K                    �?� [:��?Z           ��@G       J                    !@�ʹhrd�?           0z@H       I                    @t/*�?C            �W@������������������������       �                     0@������������������������       �        5            �S@������������������������       �        �            Pt@L       W                     @���I���?=            �[@M       R                    @�<ݚ�?             ;@N       O                    @r�q��?             2@������������������������       �        	             (@P       Q                    �?      �?             @������������������������       �                     @������������������������       �                     @S       V                    @�q�q�?             "@T       U                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @X       [                    @*�s���?+             U@Y       Z                    @nM`����?             G@������������������������       �                     =@������������������������       �                     1@������������������������       �                     C@]       �                    @*�b����?�           ��@^       i                    �?pDMM���?D           ��@_       d                     @�-ῃ�?+            �N@`       a                    @�GN�z�?             6@������������������������       �                     .@b       c                    @����X�?             @������������������������       �                     �?������������������������       ��q�q�?             @e       f                     @��Zy�?            �C@������������������������       �                     @g       h                    @     ��?             @@������������������������       �                     6@������������������������       �                     $@j                           @����-�?           ��@k       z                    �?�u��+	�?S           �@l       o                     @�q�q�?             B@m       n                    @d}h���?	             ,@������������������������       �                     @������������������������       �                     &@p       u                     @8�A�0��?             6@q       r                    �?�q�q�?             (@������������������������       �                      @s       t                    @      �?             $@������������������������       �                     @������������������������       �                     @v       y                    �?���Q��?             $@w       x                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @{       |                    @�������?=           �@������������������������       �        �            �p@}       ~                    �?Xsj�]�?�            @n@������������������������       �                      @������������������������       �        �            @m@�       �                    @x�{u��?�           |�@�       �                    �?|T����?[           ��@�       �                    @����F��?           `|@�       �                    @����X��?J            �^@������������������������       �                     ,@������������������������       �        E            @[@�       �                     @"a����?�            �t@�       �                     @j���� �?Y             a@�       �                    @ҷ{�&�?E            �Z@������������������������       �        3             T@������������������������       �                     ;@������������������������       �                     =@�       �                    @�Ha�3�?x            `h@������������������������       �        S            `a@������������������������       �        %             L@�       �                    �?�����Y�?@           P�@������������������������       �        �             n@�       �                    @&Eȧ��?�            �q@������������������������       �        -             Q@�       �                    @�8l�9��?�            �j@������������������������       �                    �E@������������������������       �        g            `e@�       �                    @��Oe� �?k           x�@�       �                    @PN���?:            @V@������������������������       �        *            �N@������������������������       �                     <@�       �                    #@�h��h�?1           ��@�       �                    �?���G�?�           x�@������������������������       �        �            �l@�       �                     @�T%��?�            �x@�       �                    @д>��C�?�            �u@�       �                    @��t����?�             j@������������������������       �        w            �f@������������������������       �                     ;@�       �                     @T�iA�?W            �a@�       �                    @z��R[�?-            �Q@������������������������       �        %            �L@������������������������       �                     *@�       �                    @����X�?*            �Q@�       �                    @�LQ�1	�?             7@������������������������       �                      @������������������������       �                     .@�       �                    @�*/�8V�?            �G@������������������������       �                     E@������������������������       �                     @������������������������       �                     G@�       �                    @��ē*�?�            pp@�       �                    @�#-���?�            �n@�       �                    @�<ݚ�?             B@������������������������       �                     <@������������������������       �                      @�       �                     @�R��ݽ?�             j@�       �                    �? �#�Ѵ�?;            �U@�       �                    %@�<ݚ�?             2@�       �                    �?X�<ݚ�?             "@������������������������       ����Q��?             @�       �                    @      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                     "@������������������������       �        .             Q@�       �                    �?��p\�?K            �^@�       �                     @@�0�!��?!            �I@�       �                    %@ �Cc}�?             <@�       �                    @�θ�?             *@�       �                    �?؇���X�?             @������������������������       �r�q��?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �        	             .@�       �                    %@��+7��?             7@�       �                    �?և���X�?             ,@������������������������       �                     @������������������������       �z�G�z�?             $@������������������������       �                     "@������������������������       �        *             R@������������������������       �                     2@�       �                    @�3��Z��?y           ��@�       �                    �?�M;q��?7            �R@������������������������       �                    �D@�       �                     @ҳ�wY;�?             A@�       �                    "@�t����?             1@������������������������       �                     @�       �                    @�q�q�?	             (@������������������������       �z�G�z�?             @������������������������       �և���X�?             @������������������������       �                     1@�       �                    �?�{�7u�?B           ��@�       �                    !@�JS���?           �{@�       �                     @�=C|F�?�            Pp@������������������������       �        @             ^@�       �                    @��|�5��?Z            �a@�       �                    @�%^�?S             `@������������������������       �                     9@�       �                     @>�Q��?C             Z@�       �                    �?ι�~��?6            �U@�       �                    @�+e�X�?             I@������������������������       �                     (@������������������������       �                     C@�       �                    @<ݚ)�?             B@�       �                    @@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@�       �                    @�eP*L��?             6@������������������������       �                     $@������������������������       �        	             (@�       �                    @X�<ݚ�?             2@������������������������       �                     $@������������������������       �                      @������������������������       �                     (@������������������������       �        t            �f@�                          !@�W(@P�?4           p@�       �                     @R��ba��?�            �s@�       �                     �?�;y�?P            �a@������������������������       �                     @�       �                    �?
�8q���?N             a@������������������������       �                     "@�       �                    �?     ��?H             `@������������������������       �                     &@�       �                    @ ���J��?C            @]@�       �                    @l��\��?             A@������������������������       �                     �?�       �                    @�FVQ&�?            �@@������������������������       �                     ?@������������������������       �                      @������������������������       �        -            �T@�       �                    �?��R���?j            �e@������������������������       �                     @                          @JF���?e            �d@                         @�q�q�?3            @T@                         @��Q��?             D@������������������������       �                     :@������������������������       �        
             ,@                         @�4F����?            �D@������������������������       �                     <@������������������������       �                     *@                         @Ї?��f�?2            @U@	      
                   �?Fmq��?!            �J@������������������������       �                     $@                         !@�%^�?            �E@                         @ �q�q�?             8@������������������������       �        	             0@                         @      �?              @������������������������       �                     �?������������������������       �                     @                         @�\��N��?             3@                         @�θ�?	             *@������������������������       �                     @������������������������       �                     $@������������������������       �                     @                         @      �?             @@������������������������       �                     (@������������������������       �                     4@������������������������       �        z            �g@�t�b�values�h,h/K ��h1��R�(KMKK��hJ�B�       8�@     ��@     `t@      D@     @k@              [@      D@              .@      [@      9@     �O@      @      0@      @      0@                      @     �G@             �F@      2@      ?@      @       @      @       @                      @      7@              ,@      .@      ,@      @      ,@      @      ,@                      @              �?              &@     ��@     >�@     �w@     �@     @l@     �@     �U@     �h@             �h@     �U@             `a@      �@     @Y@     (�@             (�@     @Y@      P@      M@      =@     �B@      =@      >@              @      =@      @      =@              <@      @      �?      @                      �?      @              5@             �E@     �A@      @      2@      @                      2@     �C@      1@     �@@      @      3@      @              @      3@              ,@              @      &@      @               @      &@              &@       @              C@     ؊@             Њ@      C@      �?      "@      �?       @      �?       @                      �?      @              =@             �b@     �w@     �S@     Pu@     �S@      0@              0@     �S@                     Pt@     @R@      C@      @      5@      @      .@              (@      @      @      @                      @      @      @      @       @      @                       @              @     �P@      1@      =@      1@      =@                      1@      C@             ��@     ��@     b�@     �|@      6@     �C@      @      1@              .@      @       @      �?              @       @      1@      6@      @              $@      6@              6@      $@             6�@     pz@     x�@      4@      8@      (@      &@      @              @      &@              *@      "@      @      @       @              @      @              @      @              @      @      �?      @      �?                      @      @             p@       @     �p@             @m@       @               @     @m@             0�@     0y@     ��@     @q@     �k@      m@     @[@      ,@              ,@     @[@              \@     `k@      L@      T@      ;@      T@              T@      ;@              =@              L@     `a@             `a@      L@             �}@     �E@      n@             �m@     �E@      Q@             `e@     �E@             �E@     `e@             ��@     �_@     �N@      <@     �N@                      <@     ��@     �X@     ��@      N@     �l@             �t@      N@      r@      N@     �f@      ;@     �f@                      ;@     �Z@     �@@     �L@      *@     �L@                      *@      I@      4@       @      .@       @                      .@      E@      @      E@                      @      G@              l@     �C@      l@      5@      <@       @      <@                       @     �h@      *@     �T@      @      ,@      @      @      @       @      @      @      �?       @              �?      �?      "@              Q@             �\@      "@      E@      "@      9@      @      $@      @      @      �?      @      �?      �?              @       @      .@              1@      @       @      @              @       @       @      "@              R@                      2@     `�@      }@      6@     �J@             �D@      6@      (@      @      (@              @      @      @      �?      @      @      @      1@             ��@     �y@     �l@     �j@     �l@     �@@      ^@              [@     �@@      X@     �@@      9@             �Q@     �@@     �O@      7@      C@      (@              (@      C@              9@      &@      *@      �?              �?      *@              (@      $@              $@      (@               @      $@              $@       @              (@                     �f@      s@     �h@      ]@     �h@      7@     �]@              @      7@     �\@      "@              ,@     �\@      &@              @     �\@      @      ?@      �?               @      ?@              ?@       @                     �T@     @W@     �S@      @             �U@     �S@      K@      ;@      :@      ,@      :@                      ,@      <@      *@      <@                      *@     �@@      J@      5@      @@      $@              &@      @@      �?      7@              0@      �?      @      �?                      @      $@      "@      $@      @              @      $@                      @      (@      4@      (@                      4@     �g@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�BX)         8                    �?.�et���?+           c�@                           @��`���?�	           0�@                           @�#Z�\�?.           x�@������������������������       �        L           ��@                           �?ދo|LL�?�           ,�@������������������������       �        ,            }@                            @������?�           �@                           !@`5)}JK�?�           8�@	       
                    @@\V�vٓ?�           (�@������������������������       �        {            �i@                           @ ��o��?           �y@                           �?��v��?�            @o@                            �?�>����?4            @T@������������������������       �                      @                           !@ �\���?2            �S@������������������������       �        ,            �Q@                            @      �?              @������������������������       �      �?             @������������������������       �      �?             @������������������������       �        f             e@������������������������       �        l            �c@������������������������       �                      @                            @ ���3�?3            }@������������������������       �                     7@                           !@��p����?"           �{@������������������������       �                   �x@                           !@�IєX�?            �I@������������������������       �                     H@������������������������       �                     @       #                     @�-�|�ʹ?d           p�@                            @���?!           �@������������������������       �        o           (�@!       "                    @��ś��?�            @q@������������������������       �        �            `o@������������������������       �                     9@$       %                    @�'�=z��?C            �X@������������������������       �                     A@&       7                    %@��&����?,            @P@'       (                    #@z�G�z�?(             N@������������������������       �                     "@)       ,                     �?������?"            �I@*       +                    @z�G�z�?             @������������������������       �      �?              @������������������������       �                     @-       .                     @�㙢�c�?             G@������������������������       �                     3@/       6                     @l��
I��?             ;@0       1                    @�㙢�c�?             7@������������������������       �                     @2       5                    @      �?
             0@3       4                     @�q�q�?             (@������������������������       ����Q��?             @������������������������       �����X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @9       :                    �?lͩ���?�           ��@������������������������       �        �           x�@;       L                    �?�j�����?�           p�@<       =                    �?��W(�!�?Q            �a@������������������������       �                     5@>       ?                    "@���*�?F             ^@������������������������       �        %            �P@@       G                    @�5��?!             K@A       D                     @p9W��S�?             C@B       C                    @D�n�3�?             3@������������������������       �                     &@������������������������       �                      @E       F                    @�S����?             3@������������������������       �                     0@������������������������       �                     @H       I                     �?     ��?
             0@������������������������       �                     @J       K                     @8�Z$���?             *@������������������������       �����X�?             @������������������������       �                     @M       �                    !@�⒱`�?�           <�@N       �                    !@��%�[H�?�           ��@O       P                    @�;,;�?<           h�@������������������������       �        [            @b@Q       r                    @l������?�           ؆@R       W                    @8����?�            �r@S       V                    @ܴD��?B            @Y@T       U                    @��x_F-�?$            �I@������������������������       �                    �D@������������������������       �                     $@������������������������       �                     I@X       Y                    �?8�A�0��?�            �h@������������������������       �                     B@Z       [                    @�E��ӭ�?f            @d@������������������������       �        $             N@\       m                     @�ʻ����?B            �Y@]       ^                    �?�c�Α�?!             M@������������������������       �                      @_       d                     �?      �?             L@`       c                    @      �?             2@a       b                    @�	j*D�?             *@������������������������       �                     "@������������������������       �                     @������������������������       �                     @e       j                    @�?�'�@�?             C@f       g                    @�nkK�?             7@������������������������       �                     @h       i                    @      �?             0@������������������������       �                     �?������������������������       �                     .@k       l                    @������?             .@������������������������       �                     @������������������������       �                     &@n       o                     @�X���?!             F@������������������������       �                     �?p       q                    @8�$�>�?             �E@������������������������       �                     <@������������������������       �                     .@s       �                     @�+$�jP�?            {@t       }                     �?@�9���?�            `l@u       |                    @>A�F<�?             C@v       w                    @l��\��?             A@������������������������       �                     �?x       {                    @�FVQ&�?            �@@y       z                    @      �?             0@������������������������       �        
             ,@������������������������       �                      @������������������������       �                     1@������������������������       �                     @~       �                    @�w��@�?~            �g@       �                    @@��8��?`             b@������������������������       �                     9@�       �                    @@��,*�?N            �]@������������������������       �        K             ]@������������������������       �                     @������������������������       �                    �F@�       �                    @,���i�?�            �i@������������������������       �        u            �f@������������������������       �                     9@�       �                    #@��H���?�           ��@������������������������       �        j             d@�       �                    @��Sݭg�?)           @}@�       �                     @fP*L��?�            @s@�       �                    @jdD{#E�?a            `b@�       �                    @     p�?W             `@�       �                    @�q�q�?             8@������������������������       �                     $@������������������������       �        
             ,@������������������������       �        G             Z@������������������������       �        
             3@�       �                    @�摋���?n             d@������������������������       �        !            �K@�       �                    @r�����?M            �Z@�       �                    @
j*D>�?             :@������������������������       �        	             $@�       �                    @     ��?             0@������������������������       �        
             &@������������������������       �                     @�       �                    @      �?6             T@������������������������       �                     ;@�       �                     @0��_��?$            �J@������������������������       �                     �?�       �                    @4��?�?#             J@������������������������       �                    �G@������������������������       �                     @�       �                     @���Q��?Z             d@�       �                    @,��I�?0            �U@�       �                     �?�%^�?            �E@������������������������       �                     ?@�       �                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                     �?�Ra����?             F@������������������������       �                     *@�       �                    @�חF�P�?             ?@�       �                    @�n_Y�K�?             *@������������������������       �      �?              @������������������������       ����Q��?             @������������������������       �        	             2@�       �                    @ox%�:�?*            @R@�       �                    @�^����?$            �M@������������������������       �        
             .@�       �                     @fP*L��?             F@������������������������       �                      @�       �                    @���H��?             E@�       �                    @�>4և��?             <@�       �                    �?�q�q�?
             .@������������������������       �                     $@������������������������       �                     @������������������������       �                     *@������������������������       �                     ,@������������������������       �                     ,@������������������������       �        �            �r@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B�       ��@     6�@     ܑ@     B�@     ��@     8�@             ��@     ��@     �}@              }@     ��@      &@     ��@       @     ��@      @     �i@             0y@      @     �n@      @     �R@      @               @     �R@      @     �Q@              @      @       @       @       @       @      e@             �c@                       @     �|@      @      7@             �{@      @     �x@              H@      @      H@                      @     @R@     L�@      9@     ��@             (�@      9@     `o@             `o@      9@              H@     �I@              A@      H@      1@      H@      (@      "@             �C@      (@      �?      @      �?      �?              @      C@       @      3@              3@       @      3@      @      @              (@      @       @      @      @       @      @       @      @                      @              @     ��@     �@     x�@             ��@     �@     �E@     �X@      5@              6@     �X@             �P@      6@      @@      &@      ;@       @      &@              &@       @              @      0@              0@      @              &@      @              @      &@       @      @       @      @             ܕ@     �y@     (�@     �y@     h�@      r@     @b@             �{@      r@     �V@      j@      $@     �V@      $@     �D@             �D@      $@                      I@     @T@     @]@      B@             �F@     @]@              N@     �F@     �L@      0@      E@       @              ,@      E@      "@      "@      "@      @      "@                      @              @      @     �@@      �?      6@              @      �?      .@      �?                      .@      @      &@      @                      &@      =@      .@      �?              <@      .@      <@                      .@      v@      T@     �e@     �K@      ?@      @      ?@      @              �?      ?@       @      ,@       @      ,@                       @      1@                      @     �a@      H@     �a@      @      9@              ]@      @      ]@                      @             �F@     �f@      9@     �f@                      9@     �@      ^@      d@             �u@      ^@     0p@     �H@     �]@      =@     �]@      $@      ,@      $@              $@      ,@              Z@                      3@     �a@      4@     �K@             �U@      4@      &@      .@              $@      &@      @      &@                      @     �R@      @      ;@              H@      @      �?             �G@      @     �G@                      @     @V@     �Q@     �B@      I@      @@      &@      ?@              �?      &@      �?                      &@      @     �C@              *@      @      :@      @       @       @      @      @       @              2@      J@      5@      J@      @      .@             �B@      @               @     �B@      @      7@      @      $@      @      $@                      @      *@              ,@                      ,@     �r@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�'         :                    �?n-����?           c�@                           @�Q���?X	           ��@                           @�
[���?           �@������������������������       �        D           ȋ@                           �?�J�{\�?�           ,�@                           !@�S�u�?S           h�@                           !@�!��b�?O           0�@������������������������       �        )            }@	       
                    @�>����?&             K@������������������������       �                     <@                           @8�Z$���?             :@                            @���Q��?	             $@                            �?���Q��?             @������������������������       �                     �?������������������������       �      �?             @                            @z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     0@������������������������       �                     @                           @�	����?           ��@������������������������       �        Z           P�@������������������������       �        %           @}@       '                     @��M�6��?B           �@                            @`1&dl�?U           Ȁ@                           @��I��?;           @������������������������       �        �            �v@                           !@��U�=��?Q            �`@������������������������       �                     1@������������������������       �        I            �\@                            @      �?             D@������������������������       �                     $@!       &                    !@�q�q�?             >@"       %                    @�LQ�1	�?             7@#       $                    @      �?              @������������������������       �                     @������������������������       �      �?             @������������������������       �        	             .@������������������������       �                     @(       +                    �?�G� �?�           @�@)       *                    @�G�z��?
             4@������������������������       �                     "@������������������������       �                     &@,       -                    @�$:b��?�           ��@������������������������       �        �            Py@.       9                    !@0aw˕��?�            �w@/       8                    @@4և���?�            �m@0       7                    @ g���B�?�            �l@1       4                     @���}<S�?=             W@2       3                    @ףp=
�?!             I@������������������������       �                    �E@������������������������       �����X�?             @5       6                    @@4և���?             E@������������������������       �                     B@������������������������       �      �?             @������������������������       �        W             a@������������������������       �                     "@������������������������       �        V             b@;       �                     @�Ϙ�.	�?�           <�@<       U                    @&��M0��?W           $�@=       T                    @Jܤm6�?�            �i@>       E                    @l�Ӑ���?n            �e@?       @                    @���� �?            �D@������������������������       �                     :@A       B                     �?������?             .@������������������������       �                      @C       D                    �?8�Z$���?             *@������������������������       �        	             &@������������������������       �                      @F       S                    !@�1��!�?P            �`@G       N                     �?�.�+��?1            �U@H       K                    @�KM�]�?             �L@I       J                    @ܷ��?��?             =@������������������������       �                     @������������������������       �                     :@L       M                    @ �Cc}�?             <@������������������������       �                     9@������������������������       �                     @O       P                    @�q�q�?             >@������������������������       �                     1@Q       R                    �?�θ�?             *@������������������������       �                     $@������������������������       �                     @������������������������       �                     G@������������������������       �                     >@V       W                    �?\=���]�?�           ��@������������������������       �        �            Pv@X       �                    @�F.< �?�           ��@Y       b                    @����n�?�           P�@Z       [                     �?�L.���?f            �c@������������������������       �                     E@\       ]                    @���Q��?N            �\@������������������������       �                     $@^       _                    @^������?F            @Z@������������������������       �                      F@`       a                    �?Nd^����?&            �N@������������������������       �                     B@������������������������       �                     9@c       d                    @ToC�g��?^           h�@������������������������       �        �            �n@e       t                    @      �?�            �s@f       g                    �?V��z4�?(             O@������������������������       �                     �?h       m                     �?�̚��?'            �N@i       j                    @      �?             >@������������������������       �                     *@k       l                    @�t����?             1@������������������������       �                     .@������������������������       �                      @n       o                    "@��a�n`�?             ?@������������������������       �                     �?p       q                    @��S�ۿ?             >@������������������������       �                     4@r       s                    @z�G�z�?             $@������������������������       �                     �?������������������������       ��<ݚ�?             "@u       v                    !@HP�s��?�            @o@������������������������       �                     $@w       x                    #@ �q�q�?�             n@������������������������       �        3             U@y       ~                    @ ��Ou��?a            �c@z       }                    �? 4^��?J            �]@{       |                     �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        G            �\@       �                    !@���"͏�?            �B@�       �                    @��H�}�?             9@�       �                     �?�n_Y�K�?             *@������������������������       �                     �?������������������������       ��q�q�?             (@�       �                    @�q�q�?	             (@������������������������       �                      @������������������������       �                     @������������������������       �                     (@������������������������       �        4            �S@�       �                     @p~i��n�?W           T�@�       �                    @��pBI�?+            @R@������������������������       �        *            �Q@������������������������       �                      @�       �                    �?^�=���?,           0�@�       �                    @d,���O�?!            �I@������������������������       �                     C@������������������������       �                     *@�       �                    @T�4��?           d�@�       �                    @��u����?j             c@�       �                    @���b��?Y             _@�       �                    @���N8�?             5@������������������������       �                     @������������������������       �                     0@�       �                    @���z�k�?I            �Y@������������������������       �        "            �G@�       �                    @����>4�?'             L@������������������������       �                     &@������������������������       �                    �F@������������������������       �                     =@�       �                    @�g+�6�?�            �@�       �                    @ �����?r           ��@������������������������       �        �            r@�       �                     @��)�1�?�           ��@�       �                    @���X��?�             l@�       �                    @x
�==Q�?~            �g@������������������������       �        +            @R@�       �                    @�����H�?S            @]@�       �                    �?x��}�?)            �K@������������������������       �        !             E@������������������������       �                     *@������������������������       �        *             O@�       �                    !@��.k���?             A@�       �                    @�n_Y�K�?             :@�       �                    �?�S����?
             3@������������������������       �                     @������������������������       �        	             0@������������������������       �                     @������������������������       �                      @�       �                    @�,_���?5            @�       �                    �?�4�����?)             O@������������������������       �                     E@������������������������       �                     4@������������������������       �                   @{@������������������������       �        /            @S@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�BP       :�@     ��@     ��@     ��@     ��@     `�@             ȋ@     ��@     �}@     �@      &@     �@      @      }@              I@      @      <@              6@      @      @      @       @      @              �?       @       @      @      �?       @               @      �?      0@                      @     P�@     @}@     P�@                     @}@     @P@      �@     �B@     @@      1@      ~@             �v@      1@     �\@      1@                     �\@      4@      4@              $@      4@      $@      4@      @      @      @      @              �?      @      .@                      @      <@     `�@      &@      "@              "@      &@              1@     �@             Py@      1@     �v@      1@     �k@       @     �k@       @      U@      @     �F@             �E@      @       @      @     �C@              B@      @      @              a@      "@                      b@     `�@     �~@     �@      q@     �]@     �U@     �]@      L@      &@      >@              :@      &@      @               @      &@       @      &@                       @     �Z@      :@     �N@      :@     �I@      @      :@      @              @      :@              9@      @      9@                      @      $@      4@              1@      $@      @      $@                      @      G@                      >@     �@     @g@     Pv@             ��@     @g@     ��@      [@      V@     @Q@      E@              G@     @Q@      $@              B@     @Q@              F@      B@      9@      B@                      9@     0�@     �C@     �n@             q@     �C@     �E@      3@              �?     �E@      2@      .@      .@              *@      .@       @      .@                       @      <@      @              �?      <@       @      4@               @       @      �?              @       @     �l@      4@              $@     �l@      $@      U@             @b@      $@     �]@      �?      @      �?              �?      @             �\@              <@      "@      0@      "@       @      @              �?       @      @       @      @       @                      @      (@                     �S@     ܑ@     �k@     �Q@       @     �Q@                       @     ��@     �k@      *@      C@              C@      *@             ��@     �f@     @X@      L@     @X@      ;@      @      0@      @                      0@      W@      &@     �G@             �F@      &@              &@     �F@                      =@     �@     �_@     �@     �H@     r@             �@     �H@     `h@      =@      f@      *@     @R@              Z@      *@      E@      *@      E@                      *@      O@              2@      0@      $@      0@      @      0@      @                      0@      @               @             �}@      4@      E@      4@      E@                      4@     @{@                     @S@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKihbh,h/K ��h1��R�(KKi��hi�B�                             @n-����?�           c�@                           �?�P[f:�?I           ��@������������������������       �        �            Ps@������������������������       �        �            �@                           �?�~@*���?�
           �@                            @@�z�'�?            �@                           �?@x�5?�?^            �@                           !@ ������?�            �o@	       
                    !@ >��@�?�            @o@������������������������       �        ~            �k@                            �?��S�ۿ?             >@������������������������       �        
             6@                           @      �?              @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �        �            @t@                           �?����|��?�            �@                           !@p/k%��?�            @t@                           !@@=��?�            �s@������������������������       �        �            �p@                           @`Ӹ����?            �F@������������������������       �                     :@                            @�KM�]�?             3@������������������������       �                     &@                           @      �?              @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        �            �w@       6                    @���)�?�           ̧@        %                    �?vw��<��?           ȉ@!       $                    @����� �?J           8�@"       #                    @��
ц��?             :@������������������������       �        	             ,@������������������������       �                     (@������������������������       �        9           �~@&       5                    �? �&�eZ�?�             s@'       (                    �?>���Rp�?#             M@������������������������       �                     ;@)       .                    @`՟�G��?             ?@*       +                     �?      �?	             0@������������������������       �                     @,       -                    @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@/       0                     �?��S���?
             .@������������������������       �                     @1       4                     @�z�G��?             $@2       3                    "@և���X�?             @������������������������       �                      @������������������������       �z�G�z�?             @������������������������       �                     @������������������������       �        �             o@7       8                    @�C�N�~�?�           Z�@������������������������       �                   �y@9       h                    @�7���?�           H�@:       ;                    �?����?�           �@������������������������       �                     @<       =                    @`�ݫ�Q�?�           ��@������������������������       �        �            Pr@>       g                    !@�C����?*           Њ@?       @                    @dP-���?!           p�@������������������������       �        	             2@A       H                     �?���.�6�?           ��@B       C                    @���|���?/            �P@������������������������       �                     >@D       E                    @�q�q�?             B@������������������������       �                     "@F       G                    �?X�<ݚ�?             ;@������������������������       �                     (@������������������������       �        	             .@I       V                    @�m(']�?�           Ї@J       K                    #@�b��fl�?b           @�@������������������������       �        �            @w@L       U                     @P���Q�?i            �f@M       N                    @�8��8��?A             [@������������������������       �                    �G@O       R                     @f>�cQ�?$            �N@P       Q                    �?0��_��?            �J@������������������������       �X�Cc�?             ,@������������������������       �                    �C@S       T                    �?      �?              @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �        (             R@W       f                     @ףp=
�?�            @j@X       Y                    �?���o��?E            �[@������������������������       �        /             R@Z       _                    @�s��:��?             C@[       \                    "@X�Cc�?	             ,@������������������������       �                     @]       ^                    @�eP*L��?             &@������������������������       �      �?             $@������������������������       �                     �?`       a                    �?      �?             8@������������������������       �                     @b       e                    @p�ݯ��?             3@c       d                    "@     ��?	             0@������������������������       �                     @������������������������       ��z�G��?             $@������������������������       �                     @������������������������       �        B             Y@������������������������       �        	             (@������������������������       �        �           x�@�t�bh�h,h/K ��h1��R�(KKiKK��hJ�B�       :�@     ��@     Ps@      �@     Ps@                      �@     Ч@     ��@     ȓ@      ,@     ��@      @      o@      @      o@       @     �k@              <@       @      6@              @       @      @              �?       @               @     @t@             ��@      $@     �s@      $@     �s@       @     �p@             �E@       @      :@              1@       @      &@              @       @      �?       @      @                       @     �w@             ؛@     ��@      s@     H�@      (@     �@      (@      ,@              ,@      (@                     �~@     @r@      ,@      F@      ,@      ;@              1@      ,@      $@      @              @      $@      �?              �?      $@              @       @              @      @      @      @      @               @      @      �?      @              o@             �@     8�@     �y@             ��@     8�@     ��@      V@              @     ��@      U@     Pr@             0�@      U@     0�@      R@              2@     0�@      K@      E@      8@      >@              (@      8@              "@      (@      .@      (@                      .@     ��@      >@     ��@      "@     @w@             `e@      "@     �X@      "@     �G@              J@      "@      H@      @      "@      @     �C@              @      @       @      @       @              R@             �g@      5@     @V@      5@      R@              1@      5@      @      "@              @      @      @      @      @              �?      (@      (@      @              @      (@      @      "@              @      @      @              @      Y@                      (@             x�@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B(          :                    �?4�L�R��?�           c�@                           @
Ic`���?B	           l�@������������������������       �                   ��@       !                    @tJ{��?&           �@                           �?��=��!�?�           ��@������������������������       �        &            |@                           !@�y��$�?�           ؐ@������������������������       �        G           ��@	                            �?�Zl�i��?n            @d@
                           �? 7���B�?"             K@                           @�KM�]�?             3@������������������������       �                     &@                           @      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                    �A@                            �?H�ՠ&��?L             [@                            @����X�?$            �H@                           @X�<ݚ�?             "@������������������������       �                     @������������������������       ��q�q�?             @                           !@      �?             D@                           @�t����?             A@������������������������       �                     .@                            @���y4F�?             3@                           @"pc�
�?	             &@������������������������       ����Q��?             @������������������������       �                     @                           @      �?              @������������������������       ����Q��?             @������������������������       �                     @������������������������       �                     @������������������������       �        (            �M@"       #                    �?(��R%��?K           ��@������������������������       �                   @{@$       +                     �?      �?;             X@%       *                     �?�<ݚ�?             "@&       )                    %@      �?              @'       (                    @����X�?             @������������������������       �      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?,       9                    !@�����?4            �U@-       .                    #@�C��2(�?/            @S@������������������������       �                     =@/       0                    @8��8���?             H@������������������������       �                     .@1       4                     @�'�`d�?            �@@2       3                    @�8��8��?             (@������������������������       �z�G�z�?             @������������������������       �                     @5       6                     @����X�?             5@������������������������       �����X�?             @7       8                    @����X�?             ,@������������������������       ����|���?             &@������������������������       �                     @������������������������       �                     $@;       �                    @F�sS�'�?�           Z�@<       u                    @�~�d�@�?+           ��@=       F                    �?PJL-S:�?V           <�@>       ?                    @�<�}���?L            @^@������������������������       �        ;            �W@@       E                     @������?             ;@A       B                    �?�q�q�?             (@������������������������       �                      @C       D                    "@�z�G��?             $@������������������������       �                     @������������������������       �      �?             @������������������������       �        	             .@G       H                    @�&����?
           X�@������������������������       �        �            �p@I       P                     �?�E���:�?c           8�@J       K                    @p���p�?D            �Y@������������������������       �                     @L       O                    !@�FVQ&�?A            �X@M       N                    @�q��/��?"            �H@������������������������       �                    �E@������������������������       �                     @������������������������       �                     I@Q       `                    @^ON��4�?            �@R       U                    @����?y           8�@S       T                    @��Sݭg�?            �C@������������������������       �                     =@������������������������       �                     $@V       W                    @      �?_            �@������������������������       �        )             P@X       Y                    �?��d��?6            ~@������������������������       �        "           �{@Z       _                     @(N:!���?            �A@[       \                    @      �?	             0@������������������������       �                     @]       ^                    "@X�<ݚ�?             "@������������������������       �                      @������������������������       �����X�?             @������������������������       �                     3@a       t                    !@Ba�x7��?�            �q@b       c                    �?�	��)��?w            �i@������������������������       �                     M@d       k                     @^H���+�?X            �b@e       f                    @������?'             Q@������������������������       �                     H@g       j                     @z�G�z�?             4@h       i                    @�����H�?             2@������������������������       �        	             0@������������������������       �                      @������������������������       �                      @l       o                    @�G�z��?1             T@m       n                    @�99lMt�?            �C@������������������������       �        	             ,@������������������������       �                     9@p       q                    �?���� �?            �D@������������������������       �                      @r       s                    @�θ�?            �C@������������������������       �                     >@������������������������       �                     "@������������������������       �        /            �R@v       {                     �?����԰?�           �@w       x                    @X�C��?G             \@������������������������       �                     .@y       z                    @DE�SA_�?@            @X@������������������������       �        <            @V@������������������������       �                      @|       �                    @�b��<3�?�           (�@}       ~                    �?�j��b�?(            �M@������������������������       �                     D@       �                     @�����?             3@������������������������       �                     @������������������������       �        
             *@�       �                    @@�[0)ʔ?f           x�@������������������������       �        �             m@�       �                    @�R�e1�?�           8�@�       �                     @ 7�+�0�?�            �@�       �                    @�O4R���?�            0w@�       �                    @ ��7��?�            �v@������������������������       �        h            �e@�       �                    !@��Μ�V�?y             h@������������������������       �                      @�       �                    �?�f]/U�?w            �g@������������������������       ��q�q�?             @������������������������       �        t            �g@�       �                    "@z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �        �            w@������������������������       �                     @������������������������       �        �            �l@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B0	       ��@     �@     ��@     ��@             ��@     ��@     ��@     ��@      }@              |@     ��@      0@     ��@             @b@      0@      J@       @      1@       @      &@              @       @               @      @             �A@             �W@      ,@     �A@      ,@      @      @      @               @      @      >@      $@      >@      @      .@              .@      @      "@       @      @       @      @              @       @      @       @      @                      @     �M@              R@     �|@             @{@      R@      8@       @      @       @      @       @      @       @       @              @              �?              �?     �Q@      1@     �Q@      @      =@             �D@      @      .@              :@      @      &@      �?      @      �?      @              .@      @      @       @      $@      @      @      @      @                      $@     �@     ؁@     �@     pu@     |�@      s@      4@     @Y@             �W@      4@      @      @      @       @              @      @              @      @      �?      .@             ,�@     `i@     �p@             ��@     `i@     @W@      $@              @     @W@      @     �E@      @     �E@                      @      I@             ��@      h@     `~@     @X@      $@      =@              =@      $@             �}@      Q@              P@     �}@      @     �{@              ?@      @      (@      @      @              @      @               @      @       @      3@              g@      X@     �[@      X@      M@              J@      X@      0@      J@              H@      0@      @      0@       @      0@                       @               @      B@      F@      9@      ,@              ,@      9@              &@      >@       @              "@      >@              >@      "@             �R@             L�@     �C@     @V@      7@              .@     @V@       @     @V@                       @     Џ@      0@     �J@      @      D@              *@      @              @      *@             (�@      $@      m@             �@      $@     �@      @     �v@      @     �v@      @     �e@             �g@      @               @     �g@      �?       @      �?     �g@              �?      @               @      �?       @     w@                      @             �l@�t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B8#                             @�w����?!           c�@                           �?�$����?�           �@������������������������       �        �            �r@������������������������       �        �           H�@       �                    @T�"n�?�
           �@                           �?�	t��ƴ?�           B�@                           @     ��?#             P@                           "@�g�y��?             ?@	       
                     �?������?             .@������������������������       �                     $@                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                            �?      �?
             0@������������������������       �                     @                            @$�q-�?	             *@������������������������       �r�q��?             @������������������������       �                     @                            �?�q�q�?            �@@������������������������       �                      @                           �?H%u��?             9@������������������������       �                     ,@                           @���!pc�?             &@������������������������       �                      @                            @�����H�?             "@������������������������       �z�G�z�?             @������������������������       �                     @       o                    @(��9N�?�           ¨@       8                    @j�y�?           �@       #                     �? �-n�?�           �@                            @0�,���?3            �P@������������������������       �                     C@!       "                    �? 	��p�?             =@������������������������       �                      @������������������������       �                     ;@$       7                    �? �Z&7v?�           ��@%       &                    !@ 5�x�?�           ��@������������������������       �        �           �@'       ,                     @`Ӹ����?9            �V@(       +                    %@�����H�?             2@)       *                    @      �?              @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     $@-       6                    %@������?-             R@.       5                    �?@9G��?            �H@/       2                     @�IєX�?             A@0       1                    @$�q-�?             *@������������������������       �                     @������������������������       �      �?              @3       4                    @���N8�?             5@������������������������       �        
             .@������������������������       �r�q��?             @������������������������       �        
             .@������������������������       �                     7@������������������������       �        �           @�@9       N                    @��2�ĺ?K           `�@:       M                     @����SS�?           �x@;       <                    �?p�C��?w            �f@������������������������       �        ,             S@=       L                    @�&=�w��?K            �Z@>       C                    @r�q��?             8@?       @                     �?�q�q�?             @������������������������       �                     �?A       B                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?D       K                    !@�����H�?             2@E       J                     �?8�Z$���?
             *@F       G                    �?�8��8��?	             (@������������������������       �                     @H       I                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        8            �T@������������������������       �        �             k@O       P                    "@z�G�z�?H            @_@������������������������       �                     @Q       V                    @@�r-��?D            �]@R       S                     �?�q�q�?             5@������������������������       �                     @T       U                     @�<ݚ�?	             2@������������������������       ��q�q�?             (@������������������������       �                     @W       h                    �?��l��?9            @X@X       c                     @������?             A@Y       b                    �?r�q��?             8@Z       [                    @�LQ�1	�?             7@������������������������       �                     @\       _                     �?r�q��?
             2@]       ^                    !@r�q��?             @������������������������       �                     @������������������������       �                     �?`       a                    !@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     �?d       e                    !@���Q��?             $@������������������������       �                     @f       g                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?i       n                     @���N8�?%            �O@j       k                    @ףp=
�?             >@������������������������       �                     5@l       m                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                    �@@p       �                    @�e j^�?�           L�@q       �                    %@0�Ђ�$�?           ��@r       u                    @�����a�?           �@s       t                    @���L��?*            �Q@������������������������       �                    �J@������������������������       �                     1@v       w                    #@@��<W��?�           ؈@������������������������       �        T           ��@x       �                     @��<b�ƥ?�            �l@y       �                    �?Pns��ޭ?Q            �`@z       {                     �?r�q��?             8@������������������������       �                     �?|                            @�㙢�c�?             7@}       ~                    @@�0�!��?	             1@������������������������       �                     @������������������������       ����!pc�?             &@�       �                    @r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �        B            @[@�       �                    @�a�O�??            @X@������������������������       �        '            �J@�       �                    �?`���i��?             F@������������������������       �ףp=
�?             $@������������������������       �                     A@������������������������       �        
             2@�       �                    @�X�C�?�             l@�       �                     @:ɨ��?            �@@�       �                    �?�\��N��?             3@������������������������       �                     @�       �                    "@����X�?             ,@������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     ,@�       �                    #@�,�q��?�            �g@�       �                    @ qP��B�?U             `@������������������������       �        @             Y@�       �                     �?ܷ��?��?             =@������������������������       �                     @������������������������       �                     :@�       �                    @Z��Yo��?-             O@������������������������       �                     >@�       �                    @     ��?             @@������������������������       �                     @�       �                    !@ȵHPS!�?             :@�       �                    �?      �?	             (@������������������������       �                     @������������������������       �                     "@������������������������       �        
             ,@������������������������       �        �           �@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B
       ��@     8�@     �r@     H�@     �r@                     H�@     0�@     (�@     0�@      a@      C@      :@      0@      .@      @      &@              $@      @      �?      @                      �?      (@      @              @      (@      �?      @      �?      @              6@      &@               @      6@      @      ,@               @      @               @       @      �?      @      �?      @             �@     �[@     ��@     �A@     �@      @     @P@       @      C@              ;@       @               @      ;@             �@      @     ��@      @     �@             �U@      @      0@       @      @       @      @              �?       @      $@             �Q@       @     �G@       @      @@       @      (@      �?      @              @      �?      4@      �?      .@              @      �?      .@              7@             @�@             �~@      =@     �x@      @     @f@      @      S@             �Y@      @      4@      @      @       @              �?      @      �?      @                      �?      0@       @      &@       @      &@      �?      @              @      �?      @                      �?              �?      @             �T@              k@              Y@      9@              @      Y@      2@      ,@      @              @      ,@      @       @      @      @             �U@      &@      :@       @      4@      @      4@      @      @              .@      @      @      �?      @                      �?      $@       @      $@                       @              �?      @      @      @              �?      @              @      �?              N@      @      ;@      @      5@              @      @      @                      @     �@@             �@      S@     X�@      D@     X�@      6@     �J@      1@     �J@                      1@     ��@      @     ��@              l@      @      `@      @      4@      @      �?              3@      @      ,@      @      @               @      @      @      �?      @               @      �?     @[@              X@      �?     �J@             �E@      �?      "@      �?      A@                      2@     �g@      B@      7@      $@      "@      $@      @              @      $@               @      @       @      ,@             �d@      :@     �_@      @      Y@              :@      @              @      :@             �C@      7@      >@              "@      7@      @              @      7@      @      "@      @                      "@              ,@             �@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�                             @R�����?           c�@                           @��l�d-�?�           �@                           �?xj�7�?Y           t�@������������������������       �                    �G@������������������������       �        :           ��@       	                    �?�?�Ʋ(�?0           X�@                           @�H�V��?�           L�@������������������������       �        �            �m@������������������������       �        C           (�@
                           �?�������?Q            ``@������������������������       �        (            �P@                           @     ��?)             P@������������������������       �                     @                            @���y4F�?$            �L@                           !@4�B��?            �B@                           @X�<ݚ�?             ;@������������������������       �        
             .@������������������������       �                     (@������������������������       �                     $@������������������������       �                     4@       :                    �?4�?�~�?	           �@       9                    !@*o��$!�?�           ,�@                           @pfc��?           |�@������������������������       �        �            �s@                           #@��k}��?L           0�@������������������������       �        �           ��@       2                     @p��%���?�            �i@                           @86��Z�?a            �c@������������������������       �                     F@       1                    @x�}b~|�?H            �\@       $                    �?�ݜ�?0            �S@        !                     �?p�ݯ��?             3@������������������������       �                      @"       #                     @�t����?             1@������������������������       �      �?              @������������������������       ��<ݚ�?             "@%       ,                     @����˵�?(            �M@&       +                     �? qP��B�?            �E@'       *                    %@ �q�q�?             8@(       )                    @z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     3@������������������������       �                     3@-       0                    %@      �?	             0@.       /                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     B@3       8                    �?@9G��?!            �H@4       5                    @�KM�]�?             3@������������������������       �                     "@6       7                    @z�G�z�?             $@������������������������       �����X�?             @������������������������       �                     @������������������������       �                     >@������������������������       �        p            �e@;       H                    �?\D�^���?�           ʢ@<       E                    @ٜSu��?.            @Q@=       >                    @Riv����?(             M@������������������������       �                     E@?       @                    "@     ��?             0@������������������������       �                     @A       B                     �?      �?	             (@������������������������       �                      @C       D                     @ףp=
�?             $@������������������������       �      �?             @������������������������       �                     @F       G                     �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@I       N                    @�y\����?�           @�@J       K                     �?~�EH,��?a            �b@������������������������       �        !            �K@L       M                    @��̅��?@            �W@������������������������       �                     B@������������������������       �        %            �M@O       P                    �?�_gX�.�?k           �@������������������������       �        �           ��@Q       �                    @�t�9�?�           h�@R       S                    @��q��?/           �@������������������������       �        �            �s@T       s                     @���d�?a           �@U       h                    @L��n��?9           �}@V       W                    �?�Q����?N            @\@������������������������       �                     @X       ]                    @|��?���?L             [@Y       \                    !@^(��I�?(            �K@Z       [                    �?�:�^���?"            �F@������������������������       �                     @������������������������       �                    �D@������������������������       �                     $@^       _                    @�#ʆA��?$            �J@������������������������       �                     8@`       a                    "@l��[B��?             =@������������������������       �                     @b       c                     �?�û��|�?             7@������������������������       �                     @d       g                    @�d�����?             3@e       f                    @��S�ۿ?             .@������������������������       �                     (@������������������������       ��q�q�?             @������������������������       �                     @i       j                    @��Ga��?�            �v@������������������������       �        /             Q@k       l                     �?��F�D�?�            �r@������������������������       �                      @m       r                    @�{Ęd�?�            pr@n       o                    #@ yqn�{?�            @r@������������������������       �        s            �f@p       q                    @ �O�H�?E            �[@������������������������       �        @             Z@������������������������       �؇���X�?             @������������������������       �                     @t       y                    @����q �?(           0~@u       x                    @�# ��?�            �w@v       w                    @��H�}�?             I@������������������������       �                     2@������������������������       �                     @@������������������������       �        �            �t@z       {                    �?�}�	���?D            �Y@������������������������       �                     D@|       �                    !@�q�q�?,            �O@}       ~                    @     ��?             @@������������������������       �                     3@       �                    @8�Z$���?             *@������������������������       �        
             &@������������������������       �                      @������������������������       �                     ?@������������������������       �        d            �c@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B0       .�@     ��@     �x@     ̡@     �G@     ��@     �G@                     ��@     �u@     ��@     �m@     (�@     �m@                     (�@      \@      3@     �P@             �F@      3@              @     �F@      (@      9@      (@      .@      (@      .@                      (@      $@              4@             �@     0�@     Ќ@     @     Ќ@     Pt@             �s@     Ќ@      (@     ��@             `h@      (@     �b@      $@      F@              Z@      $@      Q@      $@      (@      @               @      (@      @      @      @      @       @      L@      @      E@      �?      7@      �?      @      �?      �?              @      �?      3@              3@              ,@       @      �?       @      �?                       @      *@              B@             �G@       @      1@       @      "@               @       @      @       @      @              >@                     �e@     ��@     Pw@      3@      I@      "@     �H@              E@      "@      @              @      "@      @               @      "@      �?      @      �?      @              $@      �?              �?      $@             t�@     0t@     �V@     �M@     �K@              B@     �M@      B@                     �M@     �@     �p@     ��@             H�@     �p@     H�@     �Z@     �s@             ��@     �Z@     �y@     �P@      J@     �N@              @      J@      L@      ,@     �D@      @     �D@      @                     �D@      $@              C@      .@      8@              ,@      .@              @      ,@      "@              @      ,@      @      ,@      �?      (@               @      �?              @     pv@      @      Q@             0r@      @               @     0r@      @     0r@      �?     �f@             �[@      �?      Z@              @      �?              @     �{@     �C@     �v@      2@      @@      2@              2@      @@             �t@             �T@      5@      D@              E@      5@      &@      5@              3@      &@       @      &@                       @      ?@                     �c@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKwhbh,h/K ��h1��R�(KKw��hi�B         
                    @Nv.4���?           c�@                           �?0�Wd8��?n           �@������������������������       �        "           ��@       	                    @��8y��?L           Ȁ@                            �?d�nľ�?�            �v@������������������������       �                    �C@                           �?������?�            0t@������������������������       �        2             S@������������������������       �        �            �n@������������������������       �        n            �e@                            �?����I��?�
           �@                           @@����S�?'           $�@������������������������       �                     8@                           #@@���a��?           ē@������������������������       �        |           ؏@                           �?4\O�޵?�            �n@                           @�q�q��?$             H@������������������������       �                     5@                           @�5��?             ;@                            �?      �?             (@������������������������       �                      @                            @�z�G��?             $@                            @�q�q�?             "@������������������������       �      �?             @������������������������       ����Q��?             @������������������������       �                     �?                            @�r����?             .@                            �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �        x            �h@!       8                    �?h0(z��?m           ��@"       7                    @b��Z�?�           �@#       $                    #@�N�so�?�           X�@������������������������       �        >           `~@%       &                    @*eؓ���?}            �h@������������������������       �        :             W@'       *                     �?���Q��?C            @Z@(       )                    @d}h���?             ,@������������������������       �      �?             @������������������������       �                     $@+       6                    !@և���X�?=            �V@,       -                    @�J���?4            @S@������������������������       �                     ?@.       /                    @*
;&���?             G@������������������������       �                     *@0       5                    @�'�`d�?            �@@1       2                     @�q�q�?             8@������������������������       ����Q��?             $@3       4                     @d}h���?
             ,@������������������������       �r�q��?             @������������������������       �      �?              @������������������������       �                     "@������������������������       �        	             ,@������������������������       �        :           Ȍ@9       P                    @V&Y	"��?x           P�@:       ;                     �?pO��Hڮ?l           �@������������������������       �                     ,@<       E                    @���>�?e           ��@=       D                    �?$�q-�?            �C@>       A                    @؇���X�?             5@?       @                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @B       C                    �?�C��2(�?	             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     2@F       K                    @�i{�A}?G           p�@G       J                    �? ��WV�?             :@H       I                     @      �?             @������������������������       �      �?              @������������������������       �                      @������������������������       �                     6@L       O                    �? Y�5�n?7           ��@M       N                     @�8��8��?             (@������������������������       �      �?             @������������������������       �                      @������������������������       �        0           @�@Q       l                     @�;+Q��?           ��@R       k                    !@�H-���?           0z@S       V                    @D�n�3�?�            �v@T       U                    @�%����?|             h@������������������������       �        [            @b@������������������������       �        !            �G@W       X                    �?      �?i             e@������������������������       �                     @Y       Z                    @����0�?e            @d@������������������������       �                      G@[       j                    @�q3�M��?E             ]@\       e                    @����>4�?#             L@]       ^                    "@      �?             <@������������������������       �                     (@_       `                     �?     ��?
             0@������������������������       �                     @a       b                    �?�q�q�?             (@������������������������       �                      @c       d                    @�z�G��?             $@������������������������       �      �?              @������������������������       �                      @f       g                    "@؇���X�?             <@������������������������       �                     *@h       i                    @������?
             .@������������������������       �և���X�?             @������������������������       �                      @������������������������       �        "             N@������������������������       �        )             M@m       v                    !@������?�            �x@n       u                    @,;k�ɔ�?�            �t@o       p                    @ d��?�            �l@������������������������       �        q            �e@q       r                    @h�����?'             L@������������������������       �                     8@s       t                     @      �?             @@������������������������       �                      @������������������������       �                     >@������������������������       �        ?            �Y@������������������������       �        '            �P@�t�bh�h,h/K ��h1��R�(KKwKK��hJ�Bp       �@     ��@      r@     ��@             ��@      r@     �n@     �\@     �n@     �C@              S@     �n@      S@                     �n@     �e@             ֧@     ؓ@     ��@      &@      8@             ��@      &@     ؏@             `m@      &@     �B@      &@      5@              0@      &@      @      "@               @      @      @      @      @      �?      @       @      @              �?      *@       @      @       @      @                       @      @             �h@             ��@     ��@     `�@     ��@     `�@     �O@     `~@             �`@     �O@      W@              E@     �O@      @      &@      @      �?              $@     �C@      J@     �C@      C@              ?@     �C@      @      *@              :@      @      1@      @      @      @      &@      @      @      �?      @       @      "@                      ,@             Ȍ@     �@     0q@     ��@      3@              ,@     ��@      @      B@      @      2@      @       @       @       @                       @      $@      �?      $@                      �?      2@             `�@       @      9@      �?      @      �?      �?      �?       @              6@             ��@      �?      &@      �?      @      �?       @             @�@             ��@      p@     �p@      c@      j@      c@     @b@     �G@     @b@                     �G@     �O@     @Z@      @             �L@     @Z@      G@              &@     @Z@      &@     �F@      @      5@              (@      @      "@              @      @      @               @      @      @      @      �?               @      @      8@              *@      @      &@      @      @               @              N@      M@             `r@      Z@     `l@      Z@     `l@       @     �e@              K@       @      8@              >@       @               @      >@                     �Y@     �P@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B                             �?�Q����?�           c�@                           @��U��?�           ؜@                           #@�?�|�?v           ��@                           �? pƵHP�?t           ��@������������������������       �        	             (@������������������������       �        k            �@������������������������       �                     @                           �?��OI���?           �@	       
                    !@ d��?B           P@������������������������       �                   0{@                           !@"pc�
�?*            �P@                           @Xny��?'            �N@������������������������       �                     :@                           @z�G�z�?            �A@                            @�X����?             6@������������������������       �      �?              @                            @և���X�?             ,@������������������������       ����Q��?             @������������������������       �X�<ݚ�?             "@������������������������       �                     *@������������������������       �                     @������������������������       �        �           `�@                           �?�:�d�q�?c           -�@������������������������       �        r           T�@       8                    @�d�j7��?�           0�@                           �?������?�           ��@������������������������       �        ,             Q@       !                    @���n�?�           ��@                            @$����?,           �@                           �?rO(�o2�?�            �o@������������������������       �                    �J@������������������������       �        t             i@������������������������       �        �            �o@"       #                    �?�qu}+�?~            �f@������������������������       �                     @$       /                    @jه��?y            �e@%       &                    �?�z�N��?\            ``@������������������������       �        I            �Y@'       (                    @ �Cc}�?             <@������������������������       �                     �?)       .                     @�>����?             ;@*       -                    !@�r����?	             .@+       ,                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �        	             (@0       7                    @d}h���?             E@1       6                     @      �?             B@2       3                    @      �?             8@������������������������       �                     @4       5                    @���y4F�?             3@������������������������       �                     .@������������������������       �                     @������������������������       �                     (@������������������������       �                     @9       J                    �?��w��?           H�@:       ;                    "@�c�x��?6            @U@������������������������       �                     <@<       C                     @�^���U�?#            �L@=       >                    @д>��C�?             =@������������������������       �                     6@?       @                     �?����X�?             @������������������������       �                     �?A       B                    @r�q��?             @������������������������       �                     @������������������������       �      �?              @D       E                     @��>4և�?             <@������������������������       �                     @F       I                    @
;&����?             7@G       H                    @     ��?
             0@������������������������       �                     &@������������������������       �                     @������������������������       �                     @K       �                    @
�L����?�           ��@L       S                    @��;��?b           Ԡ@M       N                     �?�aZ/a��?l           ȁ@������������������������       �        0            �Q@O       P                    �?�IqB���?<           0@������������������������       �        �            �k@Q       R                    �?���=�/�?�            @q@������������������������       �        d             d@������������������������       �        E             ]@T       Y                    @�r�6z��?�           Ę@U       V                    @���܉Z�?�            �p@������������������������       �        <            �W@W       X                    �?��9
��?j            `e@������������������������       �                     D@������������������������       �        S            ``@Z       �                    !@�����?P           ��@[       \                    @XB���?F           d�@������������������������       �        �            �@]       p                    @x�L|���?           Ȃ@^       _                    @���ς̣?B           �@������������������������       �        J            �^@`       a                    #@�g<a�?�            x@������������������������       �        f             c@b       c                     �?@�R��?�             m@������������������������       �      �?             @d       e                    @�u��?�            `l@������������������������       �        P            �^@f       m                     @�q-�?@             Z@g       j                     @ȵHPS!�?!             J@h       i                    �?�KM�]�?             C@������������������������       �X�<ݚ�?             "@������������������������       �                     =@k       l                    �?؇���X�?             ,@������������������������       �z�G�z�?             $@������������������������       �                     @n       o                    �? pƵHP�?             J@������������������������       �      �?              @������������������������       �                     F@q       ~                     @���!���?=            �W@r       s                    !@H(���o�?$            �J@������������������������       �                     (@t       u                    #@D^��#��?            �D@������������������������       �                     @v       w                    �?<=�,S��?            �A@������������������������       �                     @x       }                    @d}h���?             <@y       z                     �?��
ц��?	             *@������������������������       �                     @{       |                    @���Q��?             $@������������������������       ����Q��?             @������������������������       �z�G�z�?             @������������������������       �        
             .@       �                     @��Y��]�?            �D@�       �                    �?��S�ۿ?
             .@������������������������       �                     �?������������������������       �        	             ,@������������������������       �                     :@������������������������       �        
             ,@������������������������       �        �            �l@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�BP       T�@     r�@     �@     ��@      1@      �@      (@      �@      (@                      �@      @             Ԓ@      (@     �~@      (@     0{@              K@      (@      K@      @      :@              <@      @      .@      @      @      �?       @      @      @       @      @      @      *@                      @     `�@             ��@     ��@             T�@     ��@     В@     �q@     �}@      Q@             �j@     �}@     �J@     p|@     �J@      i@     �J@                      i@             �o@      d@      3@              @      d@      (@      `@      @     �Y@              9@      @              �?      9@       @      *@       @      @       @      @                       @      @              (@             �@@      "@      ;@      "@      .@      "@              @      .@      @      .@                      @      (@              @             (�@     І@      6@     �O@              <@      6@     �A@      @      8@              6@      @       @              �?      @      �?      @              �?      �?      1@      &@      @              (@      &@      @      &@              &@      @              @             К@     ؄@     К@     `{@     �l@     0u@     �Q@              d@     0u@             �k@      d@      ]@      d@                      ]@     8�@     �X@     @l@      D@     �W@             ``@      D@              D@     ``@             ��@     �M@     ��@     �F@      �@             `�@     �F@     @      $@     �^@             pw@      $@      c@             �k@      $@      @      @     �k@      @     �^@             @X@      @      G@      @      A@      @      @      @      =@              (@       @       @       @      @             �I@      �?      @      �?      F@             �M@     �A@      3@      A@              (@      3@      6@      @              *@      6@      @              @      6@      @      @              @      @      @       @      @      @      �?              .@      D@      �?      ,@      �?              �?      ,@              :@                      ,@             �l@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�          "                    @��o���?	           c�@                           @��n��=�?�           �@                           �?ȕ��A|�?V           ��@������������������������       �                    �H@������������������������       �        :           ܔ@       !                    @��V�v�??           ��@                           �?($)Nɴ?�            y@������������������������       �        �             p@	                             @ Ϸ�~�?W             b@
                           !@�b��-8�?%            �O@                           @�w��#��?             I@                            �?���N8�?             5@������������������������       �                      @                           �?�S����?             3@������������������������       �        	             0@������������������������       �                     @                           @�f7�z�?             =@                            �?      �?              @                           @�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                            �?�ՙ/�?             5@                           @�z�G��?             $@������������������������       �                     �?                           @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @                           �?�eP*L��?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     *@������������������������       �        2            �T@������������������������       �        @           ��@#       @                    @��-%�F�?t	           ��@$       %                    �?�˘��?           ��@������������������������       �                   �|@&       '                    @��.P�?           �x@������������������������       �        F             [@(       ?                    @t|V)r�?�            �q@)       *                    �?4V��X�?^            `a@������������������������       �        	             ,@+       ,                     �?�8�Վ��?U            @_@������������������������       �                     ?@-       >                    !@��7 ���?>            �W@.       7                     @�Jhu4��?/            @R@/       0                    @`�Q��?             9@������������������������       �                     @1       4                    !@�GN�z�?             6@2       3                    �?      �?             (@������������������������       �                     @������������������������       �                     "@5       6                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @8       9                    @r�q��?             H@������������������������       �        	             (@:       ;                    !@�E��ӭ�?             B@������������������������       �                     2@<       =                    �?X�<ݚ�?
             2@������������������������       �                     $@������������������������       �                      @������������������������       �                     5@������������������������       �        ]             b@A       Z                    �?��GXT1�?V           �@B       I                     �?`bE�ė?�           L�@C       H                    !@�KM�]�?             C@D       G                    @�X�<ݺ?             B@E       F                    @�t����?
             1@������������������������       �        	             .@������������������������       �                      @������������������������       �                     3@������������������������       �                      @J       K                    #@�2����?�           ��@������������������������       �                   x�@L       Y                    �?�)���?�            �o@M       T                     @     ��?             H@N       Q                     @��2(&�?             6@O       P                    @r�q��?             @������������������������       �                     @������������������������       �                     �?R       S                    !@      �?             0@������������������������       �        
             ,@������������������������       �                      @U       V                    @�θ�?             :@������������������������       �                     ,@W       X                    @      �?             (@������������������������       ����Q��?             $@������������������������       �                      @������������������������       �        ~            �i@[       f                    @ D>!��?�           Ĝ@\       ]                    @�8���?�           ��@������������������������       �                     <@^       e                    �?��V��;�?�           ��@_       `                    "@l��
I��?             ;@������������������������       �                     @a       d                     @�����?             5@b       c                    @z�G�z�?             $@������������������������       �                     �?������������������������       ��<ݚ�?             "@������������������������       �                     &@������������������������       �        �           �@g       v                    �?���.��?�           �@h       u                    !@�{���?           �x@i       j                    @ !�8>��?�            Px@������������������������       �        �            @u@k       l                    @ \� ���?!            �H@������������������������       �                      @m       n                    #@������?            �D@������������������������       �        
             1@o       t                    @r�q��?             8@p       s                     @������?             1@q       r                     @�8��8��?             (@������������������������       �                     @������������������������       �r�q��?             @������������������������       ����Q��?             @������������������������       �                     @������������������������       �                     $@w       �                    @�M+"��?�           P�@x       y                    �?��P흹?c           (�@������������������������       �                      @z       {                    @�+��b�?a           �@������������������������       �        �            0p@|       }                    @     ��?�             r@������������������������       �        �            �m@~       �                     @z�):���?"             I@       �                    @�r����?             >@�       �                    @�IєX�?             1@�       �                     �?�����H�?             "@������������������������       �                     @�       �                    "@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                      @�       �                    "@�θ�?             *@������������������������       �                     @�       �                    @�z�G��?             $@�       �                     �?      �?              @������������������������       �                      @������������������������       �      �?             @������������������������       �                      @�       �                    @P���Q�?             4@������������������������       �                     @�       �                     @$�q-�?
             *@�       �                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        ~            �h@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�BP	       ��@     ̨@     {@     ��@     �H@     ܔ@     �H@                     ܔ@      x@     �@      x@      1@      p@              `@      1@      G@      1@     �@@      1@      0@      @               @      0@      @      0@                      @      1@      (@      @      @      @       @      @                       @               @      *@       @      @      @              �?      @       @      @                       @      @      @      @                      @      *@             �T@                     ��@     ��@     `�@      n@     �@             �|@      n@     �b@              [@      n@     �E@      X@     �E@      ,@             �T@     �E@      ?@             �I@     �E@      >@     �E@       @      1@      @              @      1@      @      "@      @                      "@       @       @       @                       @      6@      :@      (@              $@      :@              2@      $@       @      $@                       @      5@              b@             ��@     �r@     �@      *@      A@      @      A@       @      .@       @      .@                       @      3@                       @     ��@      "@     x�@             �n@      "@     �C@      "@      3@      @      @      �?      @                      �?      ,@       @      ,@                       @      4@      @      ,@              @      @      @      @       @             �i@             T�@     �q@     ��@      B@              <@     ��@       @      3@       @              @      3@       @       @       @      �?              @       @      &@             �@             �@      o@     �w@      6@     �w@      (@     @u@             �B@      (@               @     �B@      @      1@              4@      @      *@      @      &@      �?      @              @      �?       @      @      @                      $@     @�@     @l@     @�@      =@               @     @�@      ;@     0p@             Pp@      ;@     �m@              7@      ;@      @      :@      �?      0@      �?       @              @      �?      @              �?      �?       @               @      @      $@              @      @      @      @      @               @      @      @               @      3@      �?      @              (@      �?      @      �?      @                      �?      @                     �h@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKchbh,h/K ��h1��R�(KKc��hi�B�                             @V._q]��?           c�@                           �?�7ns�I�?�           ��@������������������������       �        �             t@������������������������       �        �           �@                           �?�H�++�?�
           ��@������������������������       �                   ��@       b                    @ȍm����?y           ��@                           @��S����?�           ��@	                           @�nq+N�?           4�@
                            @���}<S�?�            �l@                           �?z�G�z�?<             Y@                           @����X�?             @                           �?      �?             @������������������������       �                     �?������������������������       �                     @                            �?�q�q�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�חF�P�?6            @W@������������������������       �                    �B@                           �?���X�?!             L@������������������������       �                     0@                            �?      �?             D@                           @����X�?            �A@������������������������       �                     9@������������������������       �                     $@������������������������       �                     @������������������������       �        P            @`@������������������������       �        w           ��@        !                    !@�-��YZ�?�           4�@������������������������       �                     5@"       '                    @�S	�K��?�           ��@#       $                     �?��E��?F            �\@������������������������       �                    �@@%       &                    �?d�� z�?4            @T@������������������������       �                     7@������������������������       �        "             M@(       a                    !@��o۩f�?�           �@)       T                    @h8۝T�?�           p�@*       5                     �?�x
8|o�?W           H�@+       ,                    �?��a�n`�?             ?@������������������������       �                     @-       4                    @�����H�?             ;@.       3                    %@`2U0*��?             9@/       2                    �?��S�ۿ?             .@0       1                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                      @6       7                    @���c(�?>           P�@������������������������       �        Y           ��@8       K                    @�	�(�Z�?�            �w@9       J                    �?��RQJ��?�            �t@:       I                    %@xP�Fֺ�?5            @V@;       F                     @��[�8��?            �I@<       ?                    �?r֛w���?             ?@=       >                     @���Q��?             $@������������������������       �r�q��?             @������������������������       �      �?             @@       C                     @��s����?             5@A       B                    @���!pc�?             &@������������������������       �                     �?������������������������       ��z�G��?             $@D       E                    @ףp=
�?             $@������������������������       �                      @������������������������       �      �?              @G       H                    �?R���Q�?
             4@������������������������       �r�q��?             @������������������������       �؇���X�?             ,@������������������������       �                     C@������������������������       �        �            �m@L       M                    �?      �?             H@������������������������       �        	             0@N       Q                    @     ��?             @@O       P                     @��S�ۿ?             .@������������������������       �z�G�z�?             @������������������������       �                     $@R       S                     @�t����?             1@������������������������       ����Q��?             @������������������������       �                     (@U       V                    #@��+7��?)            @Q@������������������������       �                     @W       \                     @���!pc�?'            �P@X       Y                    �?      �?             @@������������������������       �                      @Z       [                    �?�q�q�?             8@������������������������       �                      @������������������������       �        	             0@]       `                    @�IєX�?             A@^       _                    �?Pa�	�?            �@@������������������������       �                     @@������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@������������������������       �        �            `n@�t�bh�h,h/K ��h1��R�(KKcKK��hJ�B0       6�@     ��@      t@     �@      t@                     �@     ��@     �@             ��@     ��@      w@     ��@     �_@     �@      4@     @j@      4@      T@      4@       @      @      �?      @      �?                      @      �?       @              �?      �?      �?      �?                      �?     �S@      .@     �B@             �D@      .@      0@              9@      .@      9@      $@      9@                      $@              @     @`@             ��@             ��@     �Z@              5@     ��@     �U@     �V@      7@     �@@              M@      7@              7@      M@             8�@     �O@     8�@     �C@     ��@      5@      8@      @              @      8@      @      8@      �?      ,@      �?      @      �?      @                      �?       @              $@                       @     ��@      ,@     ��@             �v@      ,@     �s@      &@     �S@      &@      D@      &@      7@       @      @      @      @      �?      �?      @      1@      @       @      @      �?              @      @      "@      �?       @              @      �?      1@      @      @      �?      (@       @      C@             �m@             �F@      @      0@              =@      @      ,@      �?      @      �?      $@              .@       @      @       @      (@             �I@      2@      @              H@      2@      0@      0@       @               @      0@       @                      0@      @@       @      @@      �?      @@                      �?              �?              8@             `n@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�                             @�<�=���?           c�@                            �?�1l�%��?u           b�@������������������������       �        <            �Z@                           �?�鞁��?9           ��@������������������������       �        �            @i@������������������������       �        �           ��@       �                    @>h���?�
           ��@       #                    �?��!�ٳ?�           ^�@	       
                     �?     ��?:             X@������������������������       �                     @                           �?jJA��v�?6            �V@������������������������       �                     @                            @0,Tg��?2             U@                           �?H�z�G�?             D@                           �?\X��t�?             7@������������������������       �                     @                           "@������?
             1@������������������������       �                     "@                           @      �?              @������������������������       ����Q��?             @������������������������       ��q�q�?             @                           @������?	             1@������������������������       �                     @                           �?�q�q�?             (@                           @X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @       "                    %@�Ra����?             F@                           @������?            �D@������������������������       �                     *@        !                    @@4և���?             <@������������������������       �                      @������������������������       �                     :@������������������������       �                     @$       9                     �?�	��7�?�           ��@%       8                     �?H�@>��?�             o@&       '                    @��L9���?�            `n@������������������������       �        D            @Y@(       /                    @R8h^��?X            �a@)       .                    �?ĭ����?O            @_@*       +                    !@0�)AU��?E            �\@������������������������       �        (             Q@,       -                    !@�nkK�?             G@������������������������       �                     F@������������������������       �                      @������������������������       �        
             &@0       1                    "@�IєX�?	             1@������������������������       �                     @2       7                    %@�C��2(�?             &@3       6                    �?�����H�?             "@4       5                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @:       =                    @��<�|�?           ��@;       <                    @��|Io��?�            �m@������������������������       �        �            @k@������������������������       �                     4@>       _                    @P��Su�?l           У@?       ^                    !@`�`~�.�?a           �@@       E                    #@@x�5?�?]            �@A       B                    @ tS==�f?�           ��@������������������������       �        $           Г@C       D                    �?�|���?s             f@������������������������       �        q            �e@������������������������       �                      @F       ]                     @X�.�d�?�            �q@G       H                    @86��Z�?n            �c@������������������������       �        +            �K@I       V                     @p���p�?C            �Y@J       M                    �?\-��p�?$             M@K       L                    �?�����H�?             B@������������������������       �և���X�?             @������������������������       �                     =@N       U                    %@"pc�
�?             6@O       P                    �?������?
             .@������������������������       �                     �?Q       T                    @����X�?	             ,@R       S                    @r�q��?             (@������������������������       �                     @������������������������       �      �?              @������������������������       �                      @������������������������       �                     @W       \                    �?`Ӹ����?            �F@X       Y                    @؇���X�?
             ,@������������������������       �      �?             @Z       [                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     ?@������������������������       �        X            �_@������������������������       �                     @`       u                    �?���]i��?           �@a       n                     @z�z�7��?+            @R@b       c                    #@�����?            �H@������������������������       �                     6@d       m                    %@��}*_��?             ;@e       j                     @`�Q��?             9@f       i                    !@      �?	             0@g       h                    @�θ�?             *@������������������������       �      �?              @������������������������       �                     @������������������������       �                     @k       l                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                      @o       p                    #@      �?             8@������������������������       �                     *@q       t                     @���!pc�?             &@r       s                    @z�G�z�?             $@������������������������       ����Q��?             @������������������������       �                     @������������������������       �                     �?v       �                    @@i�)ԙ�?�           ��@w       ~                    @@�y��?�           ��@x       }                    @ �H~�<x?�            u@y       z                    @ ��WV�?             :@������������������������       �                     3@{       |                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        �            ps@       �                    @��Μ�V�?�             x@������������������������       �        �            w@�       �                     @ҳ�wY;�?
             1@�       �                    "@      �?              @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     "@������������������������       �                     @������������������������       �        �           �@�t�b��     h�h,h/K ��h1��R�(KK�KK��hJ�Bp       ʩ@     ��@     @s@     ��@     �Z@             @i@     ��@     @i@                     ��@     b�@     �@     b�@     �_@     @Q@      ;@              @     @Q@      6@      @              O@      6@      7@      1@      $@      *@      @              @      *@              "@      @      @       @      @       @      �?      *@      @      @               @      @      @      @              @      @              @             �C@      @     �C@       @      *@              :@       @               @      :@                      @     ئ@     �X@     �j@     �A@     �j@      =@     @Y@             @\@      =@      \@      *@      \@       @      Q@              F@       @      F@                       @              &@      �?      0@              @      �?      $@      �?       @      �?      @      �?                      @              @               @              @     ,�@      P@     @k@      4@     @k@                      4@     x�@      F@     К@      3@     К@      (@     ��@       @     Г@             �e@       @     �e@                       @      q@      $@     �b@      $@     �K@             @W@      $@      I@       @      @@      @      @      @      =@              2@      @      &@      @      �?              $@      @      $@       @      @              @       @               @      @             �E@       @      (@       @      @      �?      "@      �?      "@                      �?      ?@             �_@                      @     @�@      9@      N@      *@     �C@      $@      6@              1@      $@      1@       @      $@      @      $@      @      @      @      @                      @      @       @      @                       @               @      5@      @      *@               @      @       @       @      @       @      @                      �?     `�@      (@     `�@      @      u@      �?      9@      �?      3@              @      �?      @                      �?     ps@             �w@      @     w@              &@      @       @      @               @       @      @      "@                      @             �@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�(         2                    @�'�V3��?            c�@                           �?(R��-��?�           h�@������������������������       �        f           H�@                           �?��8����?            ��@                           @2��:��?t           ��@                           @2m7a��?$           �|@������������������������       �        �            �w@������������������������       �        3            �T@	                            @��H�}�?P           h�@
                           @Nu�� �?�            �m@������������������������       �        b            @c@������������������������       �        7            �T@                           @O����?�             r@                           !@7T����?x            �g@                           �?<ݚ)�?\             b@                           @�7�yHx�?>            @Y@                           @0�� ��?,            �O@������������������������       �                     F@������������������������       �                     3@������������������������       �                     C@������������������������       �                    �E@������������������������       �                    �G@                           @�*v��??            @X@������������������������       �        ;            �V@������������������������       �                     @                           @��κc��?�            �p@                           �?P����?F            �\@������������������������       �                    �C@������������������������       �        *            �R@       )                    @0z���?f             c@       (                    @�����?;            �V@        '                     @h��@D��?,            �Q@!       $                     �?�������?             >@"       #                    @z�G�z�?             4@������������������������       �                     0@������������������������       �                     @%       &                    �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                    �D@������������������������       �                     4@*       1                     @`Jj��?+             O@+       .                     �?�r����?             >@,       -                    @$�q-�?             :@������������������������       �                     8@������������������������       �                      @/       0                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @@3       H                    @D������?�	           ^�@4       G                    @Ğ�H�w�?�           ��@5       6                     @]�����?�           ,�@������������������������       �        P           ��@7       F                    �?��Z�1f�?W           ȁ@8       C                    �?�V�ZA�?�            0p@9       :                    @X�@��l�?O            �`@������������������������       �        "            �L@;       >                    @����?-            @S@<       =                    @*
;&���?             G@������������������������       �                     @������������������������       �                    �C@?       @                    @�P�*�?             ?@������������������������       �                     (@A       B                    @�����?
             3@������������������������       �                     @������������������������       �                     *@D       E                    @K�|%��?M            @_@������������������������       �                     6@������������������������       �        ?            �Y@������������������������       �        �            `s@������������������������       �        F            �\@I       t                    �?�=�L��?�           �@J       K                    @P�*��?t            �@������������������������       �        (           �|@L       s                    !@������?L           ��@M       X                     �?�԰{��??           �@N       O                    !@�e���@�?2            @S@������������������������       �                     5@P       W                    %@�h����?#             L@Q       R                    @�Ń��̧?             E@������������������������       �                     4@S       V                    �?���7�?             6@T       U                    @�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �        	             ,@Y       Z                    @ 
N&M�?           �z@������������������������       �        b            `b@[       \                    #@����Q8�?�            �q@������������������������       �        e            �d@]       r                    %@�r����?F             ^@^       e                    �?|��"J�?.            @T@_       `                     @�������?             A@������������������������       �և���X�?             @a       d                    @�<ݚ�?             ;@b       c                     @ҳ�wY;�?	             1@������������������������       ��<ݚ�?             "@������������������������       �      �?              @������������������������       �                     $@f       k                     @��0{9�?            �G@g       j                    @      �?
             0@h       i                    @���Q��?             $@������������������������       �                     @������������������������       �և���X�?             @������������������������       �                     @l       m                     @��a�n`�?             ?@������������������������       �        	             0@n       o                    @z�G�z�?             .@������������������������       �                     @p       q                    @���!pc�?             &@������������������������       �      �?             @������������������������       �                     @������������������������       �                    �C@������������������������       �                     5@u       �                    @�������?9           H�@v                           @�˛��r�?�           p�@w       ~                    @     ��?�             n@x       }                    !@�U^����?n            �d@y       z                     �?L:�f@�?c            �b@������������������������       �                     @{       |                    �?�x�+���?_            @b@������������������������       �                     &@������������������������       �        W            �`@������������������������       �                     0@������������������������       �        /            @R@�       �                    �?,d��?O           ��@�       �                    "@��
P��?            �A@������������������������       �                     $@�       �                    @ �o_��?             9@�       �                     �?�q�q�?	             (@������������������������       �                     @�       �                     @�����H�?             "@������������������������       ��q�q�?             @������������������������       �                     @�       �                     �?�θ�?             *@������������������������       �                      @�       �                     @�C��2(�?	             &@������������������������       �z�G�z�?             @������������������������       �                     @�       �                    #@�Ar���?5           $�@�       �                    @�7X̱�?�           І@������������������������       �        �           �@�       �                    @�+e�X�?             9@������������������������       �                     @�       �                    @��2(&�?             6@������������������������       �                     3@������������������������       �                     @�       �                    @`�j~�ߵ?j           x�@������������������������       �                   �z@�       �                    �?�+$�jP�?V            �`@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�       �                    !@�h1�
U�?N            �_@�       �                    @      �?3             V@�       �                     @��Sݭg�?            �C@�       �                     �?��}*_��?             ;@�       �                    @�	j*D�?             *@������������������������       �                     @�       �                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                    @և���X�?             ,@������������������������       �                     @�       �                    @�q�q�?             "@������������������������       �      �?             @������������������������       �                     @������������������������       �                     (@�       �                     @ \� ���?            �H@�       �                    @
j*D>�?             :@�       �                     �?      �?             $@������������������������       �                     �?������������������������       �X�<ݚ�?             "@�       �                     �?      �?
             0@�       �                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @�       �                     @�nkK�?             7@�       �                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �        
             ,@������������������������       �                    �C@������������������������       �        M            �]@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B�       8�@     ��@      {@     �@             H�@      {@     ��@     �p@     @�@     �T@     �w@             �w@     �T@             �g@      u@     �T@     @c@             @c@     �T@             �Z@     �f@      Y@     �V@      Y@      F@     �L@      F@      3@      F@              F@      3@              C@             �E@                     �G@      @     �V@             �V@      @              d@     �Z@     �C@     �R@     �C@                     �R@     �^@      ?@      P@      ;@      P@      @      7@      @      0@      @      0@                      @      @      @      @                      @     �D@                      4@      M@      @      :@      @      8@       @      8@                       @       @       @       @                       @      @@             ئ@     �@     p�@      d@     p�@     �G@     ��@             P�@     �G@     �j@     �G@     @[@      9@     �L@              J@      9@     �C@      @              @     �C@              *@      2@              (@      *@      @              @      *@             �Y@      6@              6@     �Y@             `s@                     �\@     @�@     �@     �~@     P@             �|@     �~@      C@     �~@      1@      S@      �?      5@             �K@      �?     �D@      �?      4@              5@      �?       @      �?              �?       @              *@              ,@             �y@      0@     `b@             �p@      0@     �d@              Z@      0@     @P@      0@      9@      "@      @      @      5@      @      &@      @      @       @      @      @      $@              D@      @      (@      @      @      @      @              @      @      @              <@      @      0@              (@      @      @               @      @      @      @      @             �C@                      5@     ��@     �r@     ��@     �f@     @Z@     �`@      @@     �`@      0@     �`@      @              &@     �`@      &@                     �`@      0@             @R@             �@      H@      2@      1@              $@      2@      @       @      @              @       @      �?       @      �?      @              $@      @               @      $@      �?      @      �?      @             ��@      ?@     ��@      @     �@              3@      @              @      3@      @      3@                      @     ��@      9@     �z@             �[@      9@      @      @      @                      @     @Z@      6@     �P@      6@      =@      $@      1@      $@      "@      @              @      "@      �?      "@                      �?       @      @      @              @      @      @      �?              @      (@             �B@      (@      .@      &@      @      @              �?      @      @      $@      @      $@      �?      $@                      �?              @      6@      �?       @      �?       @                      �?      ,@             �C@                     �]@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�5         ,                    @�����?3           c�@                           �?�7��?�           h�@������������������������       �        z           0�@                           �?6�%���?           ��@������������������������       �        /            �U@       #                    !@z�?��?�           D�@                           @4���X"�?�           ��@                            �?f����c�?E           @@	       
                    @      �?             (@������������������������       �                     "@������������������������       �                     @                           @��f/w�?>           �~@������������������������       �        �            �w@                           �? 5x ��?A            �Z@������������������������       �                     @������������������������       �        ?             Z@                           �?|�����?�            �p@                           @Xny��?s            �f@������������������������       �                     5@������������������������       �        e            @d@                           �?�ҿf���?<            �T@������������������������       �                     9@                            @J�8���?+             M@                            �?z�G�z�?             D@                           @      �?             @������������������������       �                     @������������������������       �                     @                           @�t����?             A@                            @�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     <@!       "                    @�E��ӭ�?             2@������������������������       �        	             *@������������������������       �                     @$       +                    @��L�?�            0y@%       *                    @؝_[�3�?�            Pw@&       '                    �?�!�I�*�?y            �g@������������������������       �        9            @V@(       )                    �?Vβ���?@            @Y@������������������������       �        2             T@������������������������       �                     5@������������������������       �        s            �f@������������������������       �                     >@-       f                    @��)���?�	           ^�@.       E                    �?t�
�:��?�           �@/       >                    @"pc�
�?0            @S@0       7                     @��IF�E�?'            �P@1       2                     �?��p\�?            �D@������������������������       �                     @3       4                    @�8��8��?             B@������������������������       �                     <@5       6                    "@      �?              @������������������������       �                     @������������������������       ����Q��?             @8       9                    !@�J�4�?             9@������������������������       �        
             *@:       ;                     @�q�q�?
             (@������������������������       �                      @<       =                    @z�G�z�?             $@������������������������       �                      @������������������������       �                      @?       @                     �?���|���?	             &@������������������������       �                      @A       D                     @�<ݚ�?             "@B       C                    "@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     @F       [                    �?�Fy�^
�?�           t�@G       H                    @��c���?O           ��@������������������������       �        �            �l@I       T                    @ 4^��?�           P�@J       S                    �?@ڱ�~��?�           p�@K       L                    !@`���$��?�            �s@������������������������       �        �            �p@M       N                    @Hm_!'1�?            �H@������������������������       �                    �B@O       P                     @�q�q�?	             (@������������������������       ����Q��?             @Q       R                     @؇���X�?             @������������������������       �      �?             @������������������������       �                     @������������������������       �        �            w@U       V                     �?@4և���?             <@������������������������       ��q�q�?             @W       Z                     @`2U0*��?             9@X       Y                    @      �?              @������������������������       �                      @������������������������       �r�q��?             @������������������������       �                     1@\       ]                    @O�t8�?1           $�@������������������������       �                    �A@^       _                    @�L��D�?           ��@������������������������       �        ?           �@`       e                    @0�1�
�?�           ��@a       d                    @�qsT� �?�           l�@b       c                    @���s��?Q           ؀@������������������������       �        $            �M@������������������������       �        -            ~@������������������������       �        V            �@������������������������       �        6            �T@g       x                     �?Tm/秗�?�           ��@h       i                    @@4և���?�            @j@������������������������       �        d            @e@j       k                    @      �?             D@������������������������       �                     *@l       m                    "@X�<ݚ�?             ;@������������������������       �                     @n       w                    @�eP*L��?             6@o       p                    @p�ݯ��?             3@������������������������       �                      @q       v                    !@�t����?             1@r       s                    �?      �?
             0@������������������������       �                     @t       u                    �?���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @y       �                    @0ζ�_��?l           ��@z       }                    @��U/��?�            `u@{       |                    @؇>���?Z            @`@������������������������       �        D            �X@������������������������       �                     @@~       �                    �?��9O�?�            �j@       �                     @h�|�`�?4            �U@������������������������       �                     >@�       �                    @������?#             L@������������������������       �        	             1@�       �                    @Hث3���?            �C@������������������������       �                     4@������������������������       �                     3@�       �                    !@0,Tg��?M            �_@�       �                    @�d�����?+            @R@�       �                    �?�z�G��?             D@������������������������       �                     @�       �                     @^������?            �A@�       �                    @��.k���?             1@������������������������       �                      @������������������������       �                     "@�       �                    @r�q��?             2@������������������������       �        
             .@������������������������       �                     @�       �                     @���|���?            �@@������������������������       �                     (@�       �                    @և���X�?             5@������������������������       �                     (@������������������������       �                     "@������������������������       �        "            �J@�       �                     @�Q����?�            �@�       �                    @4��v�?�            `o@�       �                    !@؇���X�?             <@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?���7�?             6@������������������������       �                      @�       �                    @@4և���?	             ,@������������������������       �      �?             @������������������������       �                     $@�       �                    �?��j�`a�?�            �k@������������������������       �                     7@�       �                    !@p_�Q�?             i@�       �                     �?�q�q�?D             [@������������������������       �                     @�       �                    @�ԇ���?B            �Y@�       �                    @�q�����?2            �R@������������������������       �                     9@�       �                    @ �o_��?             I@������������������������       �                     ?@�       �                    @�d�����?             3@�       �                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                    #@և���X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     <@�       �                    @J� ��w�?;             W@������������������������       �        .             R@�       �                    �?      �?             4@������������������������       �                     @������������������������       �        	             .@�       �                    #@�e�����?�            Px@�       �                     @\mY@]��?�            �m@������������������������       �                     "@�       �                    !@���ei�?�            `l@�       �                     @6DSbq��?N             a@�       �                    @��.k���?>            �Y@�       �                    �?@-�_ .�?            �B@������������������������       �                      @������������������������       �                    �A@�       �                    @R=6�z�?%            @P@������������������������       �                     G@������������������������       �                     3@�       �                    @г�wY;�?             A@������������������������       �                     .@�       �                    @�}�+r��?	             3@������������������������       �                     2@������������������������       �                     �?�       �                    �?؇���X�?;            �V@�       �                    �? "��u�?             I@������������������������       �                    �G@������������������������       �                     @�       �                    @���?            �D@������������������������       �                     �?�       �                    �?R���Q�?             D@������������������������       �                     ?@������������������������       �                     "@�       �                    @������?f             c@�       �                    %@x�c/y[�?^            �`@�       �                     @���H��?]            �`@�       �                    !@     ��?             @@�       �                    �? �Cc}�?             <@������������������������       �        	             .@�       �                    �?�θ�?	             *@������������������������       �                      @�       �                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @�       �                    �?��T�u��?H            @Y@������������������������       �                     G@�       �                    @�2����?)            �K@������������������������       �                     @�       �                    @     ��?#             H@�       �                    �?�c�Α�?             =@�       �                    �?z�G�z�?             $@�       �                    !@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    @�����?             3@������������������������       �                     @������������������������       �        
             *@�       �                    �?�}�+r��?             3@�       �                    !@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@������������������������       �                     �?������������������������       �                     3@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�BP       ��@     <�@     �|@     Ԡ@             0�@     �|@     ��@     �U@             0w@     ��@      t@     �{@     @\@     0x@      "@      @      "@                      @      Z@      x@             �w@      Z@      @              @      Z@             �i@     �M@     @d@      5@              5@     @d@             �F@      C@      9@              4@      C@      @     �@@      @      @      @                      @      @      >@      @       @               @      @                      <@      *@      @      *@                      @     �I@      v@      5@      v@      5@      e@             @V@      5@      T@              T@      5@                     �f@      >@             ��@     ��@     T�@     �}@      ,@     �O@      @     �M@      @      C@              @      @     �@@              <@      @      @              @      @       @      @      5@              *@      @       @       @               @       @               @       @              @      @               @      @       @      @       @              �?      @      �?      @             8�@     �y@      �@     �m@             �l@      �@      @     P�@      @     �s@      @     �p@             �F@      @     �B@               @      @       @      @      @      �?      @      �?      @             w@              :@       @       @      �?      8@      �?      @      �?       @              @      �?      1@             `�@      f@             �A@     `�@     �a@     �@              �@     �a@      �@     �M@      ~@     �M@             �M@      ~@              �@                     �T@     ��@     p}@     `h@      .@     @e@              9@      .@      *@              (@      .@              @      (@      $@      (@      @               @      (@      @      (@      @      @              @      @      @                      @              �?              @     p�@     �|@      n@     �Y@     �X@      @@     �X@                      @@     �a@     �Q@     �H@     �B@      >@              3@     �B@              1@      3@      4@              4@      3@             @W@     �@@      D@     �@@      <@      (@      @              7@      (@       @      "@       @                      "@      .@      @      .@                      @      (@      5@              (@      (@      "@      (@                      "@     �J@             �q@      v@     �X@      c@      8@      @      @      @      @                      @      5@      �?       @              *@      �?      @      �?      $@             �R@     �b@      7@             �I@     �b@      B@      R@              @      B@     �P@      B@     �C@              9@      B@      ,@      ?@              @      ,@      �?      &@      �?                      &@      @      @       @               @      @       @                      @              <@      .@     @S@              R@      .@      @              @      .@             �g@      i@     �Q@     �d@      "@              O@     �d@     �H@     �U@      H@      K@       @     �A@       @                     �A@      G@      3@      G@                      3@      �?     �@@              .@      �?      2@              2@      �?              *@     �S@      @     �G@             �G@      @              $@      ?@      �?              "@      ?@              ?@      "@             @]@      B@     @]@      1@     @]@      0@      9@      @      9@      @      .@              $@      @               @      $@      �?      $@                      �?              @      W@      "@      G@              G@      "@      @             �C@      "@      5@       @       @       @       @       @       @                       @      @              *@      @              @      *@              2@      �?       @      �?       @                      �?      0@                      �?              3@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KKɅ�hi�B�+         4                    �?䀂!���?            c�@       #                    !@~�_���?�           ��@       "                    �?�������?           h�@                           @
t1���?8           x�@                            �?���I���?�            �v@������������������������       �        
             3@       
                    @6��(��?�            `u@       	                    @z���A�?�             n@������������������������       �        �            `g@������������������������       �                     K@                           @�#l��?A            @Y@                           @�e����?            �C@������������������������       �                     (@                           @�5��?             ;@������������������������       �        	             0@������������������������       �        	             &@������������������������       �        )             O@                           @�e5��o�?I           0�@������������������������       �        W            �b@                            �?��T��?�            w@                           !@���7�?             6@������������������������       �                     "@                           @$�q-�?             *@������������������������       �                     @                           @r�q��?             @������������������������       �                     �?������������������������       �                     @                           !@��|�?�w?�            �u@������������������������       �        �            @s@       !                     @ ���J��?            �C@                            @      �?              @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     ?@������������������������       �        �           X�@$       1                    !@���.�6�?�            @q@%       &                    @��}����?�            �p@������������������������       �        f             e@'       .                     @ ���3�??            �X@(       )                    @>a�����?            �I@������������������������       �                     @*       +                    �?dP-���?            �G@������������������������       �                     @,       -                    @`���i��?             F@������������������������       �                    �E@������������������������       �                     �?/       0                    �?8��8���?              H@������������������������       �                    �E@������������������������       �                     @2       3                     @      �?              @������������������������       �                     @������������������������       �                     @5       �                    @ƫ�A'��?U           ��@6       A                    @:�?���?�           J�@7       :                    @�P���R�?           <�@8       9                    �?�i��h��?\           ��@������������������������       �                     E@������������������������       �        A           ��@;       <                    �?HP�s��?�            0q@������������������������       �        3            @W@=       >                    �?Ĝ�oV4�?s            �f@������������������������       �        J            �\@?       @                    @�!���?)             Q@������������������������       �                     G@������������������������       �                     6@B       O                    @@�@K��?�           ��@C       D                    @�ٹ��?�           �@������������������������       �        t            �f@E       N                    @��vK�ݨ?N           P�@F       M                    �?�c釠�?�            �n@G       H                     @t�G����?n            �e@������������������������       �        @             Z@I       L                    @�����?.             Q@J       K                    @4և����?%             L@������������������������       �        	             *@������������������������       �                    �E@������������������������       �        	             (@������������������������       �        *            �R@������������������������       �        �            @q@P       y                    !@�!�*`M�?�           T�@Q       x                    @�����?}           ��@R       g                    �?���YU�?s           0�@S       ^                    @ �=����?�            q@T       [                    @���c���?C             Z@U       Z                    @�n���?.             R@V       W                     @�����H�?            �F@������������������������       �                     3@X       Y                    @���B���?             :@������������������������       �                     @������������������������       �                     5@������������������������       �                     ;@\       ]                    @     ��?             @@������������������������       �                     "@������������������������       �                     7@_       b                     @(.�`(�?h             e@`       a                    @����?1            �U@������������������������       �        -             T@������������������������       �                     @c       d                    @������?7            �T@������������������������       �                     D@e       f                    !@�����?             E@������������������������       �                     @������������������������       �                     C@h       s                     @ �#���?�            Ps@i       r                    @R�}e�.�?d            �c@j       k                    @؇���X�?            �H@������������������������       �                     C@l       q                    @���|���?	             &@m       p                    !@�q�q�?             @n       o                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        E            �Z@t       w                    @d=0��?d             c@u       v                    �?����0�?!             K@������������������������       �                     3@������������������������       �                    �A@������������������������       �        C            �X@������������������������       �        
             .@z       �                    @��Q���?S            �@{       �                    @և���X�?p            �e@|       }                     �?@w��_m�?S            �_@������������������������       �                     ,@~                           �?��(�?L            @\@������������������������       �        
             *@������������������������       �        B             Y@������������������������       �                     H@�       �                    %@`�|+��?�           ��@�       �                     �?Dk�-,��?�           0�@�       �                     �?8^s]e�?'             M@�       �                    �?������?%             K@������������������������       �                     @�       �                    @��[�8��?"            �I@������������������������       �                     $@�       �                    �?���� �?            �D@������������������������       �                     �?�       �                    @      �?             D@������������������������       �                     :@�       �                    @����X�?	             ,@�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?��u�s�?�           `�@�       �                    @��M9�U�?C            �[@������������������������       �        	             *@�       �                    @�q��/��?:            �X@������������������������       �                    �@@�       �                     @�����D�?'            @P@�       �                     @�����?            �H@�       �                    !@     ��?             @@�       �                    @ 	��p�?             =@�       �                    @�r����?             .@������������������������       �                     @������������������������       �      �?              @������������������������       �                     ,@������������������������       �                     @�       �                    @�t����?
             1@�       �                    @$�q-�?             *@������������������������       �                     @������������������������       �؇���X�?             @������������������������       �                     @�       �                    #@      �?             0@������������������������       �                     �?�       �                    @�r����?
             .@������������������������       �                     @�       �                    @z�G�z�?             $@������������������������       ����Q��?             @������������������������       �                     @�       �                    @��U�i:�?M           �@�       �                    @`Ӹ����?8            �V@������������������������       �                     6@�       �                     @�IєX�?+             Q@�       �                    @؇���X�?             <@�       �                    �?$�q-�?             :@������������������������       ��q�q�?             @�       �                    @�nkK�?             7@������������������������       �                     0@������������������������       �؇���X�?             @������������������������       �                      @������������������������       �                     D@�       �                    #@�!�	��?           0|@������������������������       �        m            `f@�       �                    @�IєX�?�             q@������������������������       �                    �J@�       �                     @��n5V�?�            `k@�       �                    @(2��R�?H            �]@�       �                    �? ѯ��?B            �Z@������������������������       ��q�q�?             "@������������������������       �        =            �X@�       �                    @�C��2(�?             &@������������������������       �r�q��?             @������������������������       �                     @������������������������       �        A            @Y@�       �                    @�sly47�?,            �R@������������������������       �                     J@������������������������       �                     7@������������������������       �        �           @�@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B�       p�@     V�@     (�@      �@     ��@      v@     h�@      v@     �c@     `i@      3@             `a@     `i@      K@     `g@             `g@      K@             @U@      0@      7@      0@      (@              &@      0@              0@      &@              O@             �v@     �b@             �b@     �v@       @      5@      �?      "@              (@      �?      @              @      �?              �?      @             �u@      �?     @s@              C@      �?      @      �?      @               @      �?      ?@             X�@              2@      p@      *@     �o@              e@      *@     �U@       @     �E@      @              @     �E@      @              �?     �E@             �E@      �?              @     �E@             �E@      @              @      @              @      @             \�@     ��@     \�@     ܕ@     pr@     @�@      E@     ��@      E@                     ��@     �o@      6@     @W@              d@      6@     �\@              G@      6@      G@                      6@     �@     �|@     ��@      *@     �f@             �@      *@      m@      *@     �c@      *@      Z@             �K@      *@     �E@      *@              *@     �E@              (@             �R@             @q@             L�@      |@     �t@     �p@     �t@      o@     @Y@     �e@     �V@      ,@     �P@      @      D@      @      3@              5@      @              @      5@              ;@              7@      "@              "@      7@              &@     �c@      @      T@              T@      @              @     �S@              D@      @      C@      @                      C@      m@     @S@     �\@      E@      @      E@              C@      @      @       @      @      �?      @      �?                      @      �?              @             �Z@             �]@     �A@      3@     �A@      3@                     �A@     �X@                      .@     0�@     @g@     �R@      Y@      ;@      Y@      ,@              *@      Y@      *@                      Y@      H@             ؅@     �U@     8�@     �O@      D@      2@      D@      ,@              @      D@      &@      $@              >@      &@              �?      >@      $@      :@              @      $@      @      @      @                      @              @              @     ��@     �F@     �U@      9@              *@     �U@      (@     �@@             �J@      (@     �C@      $@      ;@      @      ;@       @      *@       @      @              @       @      ,@                      @      (@      @      (@      �?      @              @      �?              @      ,@       @      �?              *@       @      @               @       @      @       @      @             H�@      4@     �U@      @      6@              P@      @      8@      @      8@       @       @      �?      6@      �?      0@              @      �?               @      D@             0{@      0@     `f@              p@      0@     �J@             `i@      0@     �Y@      0@     @Y@      @      @      @     �X@              �?      $@      �?      @              @     @Y@              J@      7@      J@                      7@             @�@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B('         ,                    @ny͈0��?           c�@                           �?"�����?�           ؤ@������������������������       �        z           @�@                           �?�|��NJ�?           p�@       
                    @����
�?a           ��@       	                    !@(=��?�?�           ȃ@                           @�'�ſ:�?!            }@������������������������       �        �            �h@������������������������       �        �            �p@������������������������       �        j             e@                           @��.N"Ҭ?�            �u@������������������������       �        a            �d@                           @����a�?u            `f@������������������������       �        o             e@������������������������       �                     $@                           @��Q�2_�?�            �p@                           �?���vq�?E            �Z@������������������������       �                    �@@������������������������       �        .            @R@       +                    !@     ��?h             d@                           @���!pc�?H            �[@                            �?�Q����?             D@������������������������       �                      @                           �?     ��?             @@������������������������       �                     &@������������������������       �                     5@       $                     �?������?,            �Q@                           @      �?             0@������������������������       �                     @       !                    @���!pc�?	             &@                            @      �?             @������������������������       �                      @������������������������       �                      @"       #                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?%       &                    �?@3����?              K@������������������������       �                    �C@'       (                    @��S�ۿ?             .@������������������������       �                     @)       *                     @      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      I@-       N                    @<4w�I��?}	           �@.       3                    �?��$�?��?           T�@/       0                     @0*��ɾ?4            @������������������������       �        �            0r@1       2                    @�n����?�            �i@������������������������       �                     @@������������������������       �        n            �e@4       E                    @ �R[u�?�           �@5       6                     �?�R�G�?P            @_@������������������������       �                    �@@7       8                     @
;&����?<             W@������������������������       �                     ;@9       :                    @@i��M��?)            @P@������������������������       �                     (@;       @                    @�iʫ{�?"            �J@<       ?                    !@���!pc�?             6@=       >                    @���Q��?             .@������������������������       �                     "@������������������������       �                     @������������������������       �                     @A       D                    !@��a�n`�?             ?@B       C                    @�S����?
             3@������������������������       �                     0@������������������������       �                     @������������������������       �                     (@F       G                    @(M�׈�?           0�@������������������������       �        �            p@H       I                    �?����n�?�            Pv@������������������������       �        .            @R@J       K                     �?�d�!۵�?�            �q@������������������������       �        !            �I@L       M                    @l��z?��?�             m@������������������������       �        o            `f@������������������������       �        &             K@O       R                    @pȬM���?z           D�@P       Q                    �?u����?�           h�@������������������������       �        O             _@������������������������       �        f           ��@S       �                    @�ZĄ��?�           ԝ@T       a                    �?0y�^E�?�           <�@U       V                    @Nd^����?)            �N@������������������������       �                     "@W       X                     �?�	j*D�?#             J@������������������������       �                     $@Y       Z                    "@؇���X�?             E@������������������������       �                     @[       \                    �?�?�|�?            �B@������������������������       �                     2@]       `                     @�}�+r��?             3@^       _                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@b       m                    @��8�$>�?Y           H�@c       l                    @x�ۈp�?d            `e@d       g                     @\X��t�?             G@e       f                    @@4և���?             ,@������������������������       �        
             *@������������������������       �                     �?h       i                     @     ��?             @@������������������������       �                     $@j       k                    @8�A�0��?             6@������������������������       �        	             *@������������������������       �                     "@������������������������       �        F            @_@n       �                    !@C��X�?�           ��@o       �                    �?��S�#�?�           p�@p       �                    �?`>:�7�?�           ��@q       x                     �?���q��?{            �g@r       s                    @ �Cc}�?             <@������������������������       �        	             *@t       u                    !@z�G�z�?             .@������������������������       �                     @v       w                    @      �?              @������������������������       �                     @������������������������       �                     @y       z                    @������?g            `d@������������������������       �        )             N@{       �                    @�]��?>            �Y@|       �                     @$�q-�?             J@}       �                     @Pa�	�?            �@@~                           !@h�����?             <@������������������������       �                     9@������������������������       ��q�q�?             @������������������������       �                     @�       �                    !@�S����?             3@������������������������       �        
             .@������������������������       �      �?             @������������������������       �                    �I@������������������������       �        F           �@�       �                     �?((8��e�?*           ��@�       �                    @�GN�z�?'            �P@�       �                    �?�C��2(�?"            �K@������������������������       �                     I@������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    #@����ۧ?           ��@�       �                     @ �>#b�?#           @|@�       �                    @ �+�^}�?�            �m@������������������������       �        V            �`@�       �                    !@��9J���?C             Z@������������������������       �                     @������������������������       �        @            @Y@������������������������       �        �            �j@�       �                    @ �#�Ѵ�?�            �u@�       �                    �?㺦���?9            @W@������������������������       �                    �C@�       �                     @H�ՠ&��?             K@�       �                    @R�}e�.�?             :@�       �                    @��2(&�?	             6@������������������������       �                     ,@������������������������       �      �?              @������������������������       �                     @������������������������       �                     <@�       �                    @�"�<F��?�            `o@�       �                    �?�� r/E�?�            �n@�       �                    @"pc�
�?             6@�       �                     @����X�?             ,@�       �                     @z�G�z�?             $@������������������������       �      �?             @������������������������       �r�q��?             @������������������������       �      �?             @������������������������       �                      @�       �                    @ >��
�?�             l@������������������������       �        �            �i@�       �                     @�����H�?             2@������������������������       ��<ݚ�?             "@������������������������       �                     "@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             &@������������������������       �        C            �Y@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B0       d�@     b�@     �{@     f�@             @�@     �{@     �@     `q@     ��@     �p@     �v@     �p@     �h@             �h@     �p@                      e@      $@     �t@             �d@      $@      e@              e@      $@             `d@     �Y@     �@@     @R@     �@@                     @R@     @`@      >@      T@      >@      3@      5@       @              &@      5@      &@                      5@     �N@      "@       @       @              @       @      @       @       @       @                       @      @      �?      @                      �?     �J@      �?     �C@              ,@      �?      @              @      �?              �?      @              I@             �@     ��@     <�@     �`@      }@      @@     0r@             �e@      @@              @@     �e@             �@     �Y@     @S@      H@     �@@              F@      H@              ;@      F@      5@              (@      F@      "@      0@      @      "@      @      "@                      @      @              <@      @      0@      @      0@                      @      (@             ��@      K@     p@             �r@      K@     @R@             �l@      K@     �I@             `f@      K@     `f@                      K@     ��@     ��@      _@     ��@      _@                     ��@     ��@     �h@     ��@     @X@      B@      9@              "@      B@      0@              $@      B@      @              @      B@      �?      2@              2@      �?      @      �?      @                      �?      ,@             (�@      R@     �b@      4@      :@      4@      *@      �?      *@                      �?      *@      3@              $@      *@      "@      *@                      "@     @_@             ̗@      J@     ̗@     �D@     ��@      @      g@      @      9@      @      *@              (@      @      @              @      @              @      @             �c@      @      N@             �X@      @      H@      @      @@      �?      ;@      �?      9@               @      �?      @              0@      @      .@              �?      @     �I@             �@             ��@      A@     �I@      .@      I@      @      I@                      @      �?      $@      �?                      $@     H�@      3@     |@      @     `m@      @     �`@             @Y@      @              @     @Y@             �j@             �t@      0@     �U@      @     �C@             �G@      @      3@      @      3@      @      ,@              @      @              @      <@             @n@      "@      n@      @      2@      @      $@      @       @       @      @      �?      @      �?       @       @       @             �k@       @     �i@              0@       @      @       @      "@              �?      @      �?                      @              &@             �Y@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKwhbh,h/K ��h1��R�(KKw��hi�B                             @KH{��?�           c�@                           @����?E           ��@                           @��5�L�?+           X�@������������������������       �        �            �@                           �?@��_;�?=            @������������������������       �        ,           P}@������������������������       �                     =@       	                     �?
3j���?           (�@������������������������       �        <            @V@
                           �?��U<�q�?�           `�@                           �?,N�_� �?�            �r@������������������������       �        �            @q@������������������������       �                     4@                           �?�G�����?+           @~@������������������������       �        Z            @b@������������������������       �        �             u@                           �?�9�gG�?�
           �@������������������������       �        D           ��@       .                    @ �$����?r           ��@       )                    �?0eg���?�           ̖@       &                    �?Vβ���??            @Y@                           @�MWl��?#            �L@                           �?�������?             A@������������������������       �        	             0@                           "@      �?             2@������������������������       �                     @                            @      �?             (@                            �?      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                      @        !                    �?�㙢�c�?             7@������������������������       �                     *@"       #                    "@���Q��?             $@������������������������       �                     @$       %                     �?؇���X�?             @������������������������       �                     �?������������������������       �                     @'       (                    @"pc�
�?             F@������������������������       �                      @������������������������       �                     B@*       -                    %@�a�O�?\           8�@+       ,                    @��]-@~?W           �@������������������������       �                     @������������������������       �        S            �@������������������������       �                     "@/       V                    @4��ƹ��?�           ��@0       U                    @L�����?�           L�@1       <                    @��v��?�           @�@2       ;                    %@؇���X�?$             L@3       4                    !@$�q-�?!             J@������������������������       �                     C@5       :                     @����X�?
             ,@6       9                     @���Q��?             $@7       8                    �?      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @=       T                    �?P����?^           ��@>       ?                    !@�&=�w��?           �z@������������������������       �        �            �s@@       O                     @f1r��g�?>            �Z@A       F                    �?ףp=
�?/             T@B       C                     �?X�<ݚ�?	             "@������������������������       �                      @D       E                     @����X�?             @������������������������       ����Q��?             @������������������������       �                      @G       N                    %@����Q8�?&            �Q@H       M                     @���y4F�?
             3@I       J                    @����X�?             ,@������������������������       �                     @K       L                     �?X�<ݚ�?             "@������������������������       �      �?             @������������������������       ����Q��?             @������������������������       �                     @������������������������       �                     J@P       S                    %@�	j*D�?             :@Q       R                    �?��S���?             .@������������������������       �                     @������������������������       ����|���?             &@������������������������       �                     &@������������������������       �        N           @�@������������������������       �        B            �Z@W       ^                    �?���l�?           ��@X       Y                    !@����?s             f@������������������������       �        b            �b@Z       [                    @д>��C�?             =@������������������������       �                      @\       ]                    !@���N8�?             5@������������������������       �        
             0@������������������������       �                     @_       v                    @Zsfi��?�           ��@`       a                    @�Ra����?f           ��@������������������������       �        �             p@b       g                    �?���?�            �s@c       d                    @Lő����?�            `j@������������������������       �        _            @b@e       f                    !@��&����?(            @P@������������������������       �                     H@������������������������       �        
             1@h       i                    �?�	��)��?>            �Y@������������������������       �                     @j       u                     @X�<ݚ�?<            �X@k       l                    �?d}h���?$             L@������������������������       �                     @m       n                    "@ i���t�?            �H@������������������������       �                     @@o       t                    @�t����?             1@p       q                     �?      �?	             $@������������������������       �                      @r       s                    @      �?              @������������������������       �      �?             @������������������������       �      �?             @������������������������       �                     @������������������������       �                    �E@������������������������       �        :            �X@�t�b��      h�h,h/K ��h1��R�(KKwKK��hJ�Bp       F�@     ��@     �q@     |�@      =@     �@              �@      =@     P}@             P}@      =@             �o@     0�@     @V@             �d@     0�@      4@     @q@             @q@      4@             @b@      u@     @b@                      u@     �@     ��@             ��@     �@     �t@     @�@     �A@      T@      5@      F@      *@      9@      "@      0@              "@      "@              @      "@      @      �?      @               @      �?      �?       @              3@      @      *@              @      @              @      @      �?              �?      @              B@       @               @      B@              �@      ,@      �@      @              @      �@                      "@     ܙ@     �r@     ��@     ``@     ��@      8@      H@       @      H@      @      C@              $@      @      @      @      @       @               @      @                       @      @                      @      �@      0@     �y@      0@     �s@             �V@      0@      R@       @      @      @               @      @       @      @       @       @             �P@      @      .@      @      $@      @      @              @      @       @       @      @       @      @              J@              2@       @      @       @              @      @      @      &@             @�@                     �Z@     8�@      e@     �e@      @     �b@              8@      @       @              0@      @      0@                      @     �@     �d@     �@     @P@      p@              o@     @P@     @h@      1@     @b@              H@      1@      H@                      1@     �K@      H@              @     �K@      F@      (@      F@      @              @      F@              @@      @      (@      @      @               @      @      @       @       @      @      �?              @     �E@                     �X@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B$         B                    �?4��1��?�           c�@                           @Z��:��?!	           �@������������������������       �                   �@       A                    @��0U��?           ȟ@       $                    @�8���+�?�           ��@       #                    �? mm�U�?�           ��@                            @0����?R           ��@                           !@@A��q�?�            �p@	                            �?�\5ݓˎ?�            �p@
                           !@�(\����?             D@������������������������       �                     6@                           @�X�<ݺ?	             2@                           @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@                           @����>4�?�             l@                           !@���=��?g            �b@������������������������       �        Y            �`@                           @      �?             0@������������������������       �                      @                            @      �?              @������������������������       �      �?             @������������������������       �                     @������������������������       �        *            �R@������������������������       �                     @                           !@����$�?�            �p@������������������������       �        �            �m@       "                    !@ȵHPS!�?             :@                           @ �q�q�?             8@������������������������       �                     (@        !                    @�8��8��?             (@������������������������       �r�q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        O           X�@%       ,                     �?�3Ea�$�?>             W@&       +                     �?X�<ݚ�?             "@'       *                    %@      �?              @(       )                    @����X�?             @������������������������       �r�q��?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?-       .                    #@4�{Y���?9            �T@������������������������       �                     ?@/       @                    %@R�}e�.�?"             J@0       7                     @d,���O�?!            �I@1       6                    !@�LQ�1	�?             7@2       3                    @�C��2(�?             6@������������������������       �                     $@4       5                    @r�q��?	             (@������������������������       �����X�?             @������������������������       �                     @������������������������       �                     �?8       ?                    @X�Cc�?             <@9       :                    @"pc�
�?             6@������������������������       �                      @;       >                    @����X�?
             ,@<       =                     @�	j*D�?	             *@������������������������       �      �?              @������������������������       ����Q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        5           ��@C       �                    @b�z�47�?�           ԥ@D       S                    �?����%��?I           �@E       F                    �?4�B��?Z            �b@������������������������       �                     6@G       H                    @Z���c��?O            �_@������������������������       �        1            �S@I       R                     @r�q��?             H@J       K                    "@¦	^_�?             ?@������������������������       �        	             ,@L       O                    @��.k���?             1@M       N                     �?X�<ݚ�?             "@������������������������       �                      @������������������������       �����X�?             @P       Q                     �?      �?              @������������������������       �                     �?������������������������       �և���X�?             @������������������������       �        
             1@T       _                    @`���Ֆ�?�           �@U       X                    @�	�{��?            ��@V       W                    @4���C�?)            �P@������������������������       �                     <@������������������������       �                     C@Y       ^                    @�Ը�p�?�           ��@Z       [                    �?�jFc�N�?�           ��@������������������������       �        �           8�@\       ]                    @��.k���?1            @U@������������������������       �                    �F@������������������������       �                     D@������������������������       �                   (�@`       �                    !@,��v4v�?�           ��@a       �                     @�����m�?           Py@b       o                    @��`h�e�?�            `k@c       d                     �?D�n�3�?             C@������������������������       �        	             ,@e       j                    @�q�q�?             8@f       g                    �?����X�?	             ,@������������������������       �                     @h       i                    "@���|���?             &@������������������������       �                      @������������������������       ��<ݚ�?             "@k       n                    "@���Q��?             $@l       m                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �z�G�z�?             @p                            �?T�<���?x            �f@q       r                    �?4��Q���?K            @\@������������������������       �                     �?s       v                    @�X�C�?J             \@t       u                    @z�G�z�?             >@������������������������       �                     8@������������������������       �                     @w       |                    @ĴF���?7            �T@x       y                    @؇���X�?             E@������������������������       �                     6@z       {                    @�z�G��?             4@������������������������       �                     ,@������������������������       �                     @}       ~                    @�(\����?             D@������������������������       �                    �C@������������������������       �                     �?�       �                    �?��M���?-             Q@������������������������       �                     @�       �                    @`��:�?(            �N@������������������������       �                     .@�       �                    @��+7��?             G@�       �                    @�z�G��?             D@�       �                    �?H%u��?             9@������������������������       �                     @������������������������       �                     6@�       �                    @���Q��?
             .@������������������������       �                     "@������������������������       �                     @������������������������       �                     @�       �                    @t�7��?{            @g@�       �                    @�8�ͻ��?P             _@������������������������       �                     0@�       �                    @<ݚ)�?H             [@�       �                    @�q�q�?             8@������������������������       �                     $@������������������������       �                     ,@�       �                    �?�/,Tg�?:             U@������������������������       �                     @�       �                    @����?4            �S@������������������������       �                    �A@�       �                    !@�+��<��?            �E@�       �                    �?�q�q�?             5@������������������������       �                     @�       �                    @��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?�       �                    �?�GN�z�?             6@������������������������       �                     $@�       �                    @�q�q�?	             (@������������������������       �                     @������������������������       �                     @������������������������       �        +             O@������������������������       �        �            �s@������������������������       �        �            �k@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�BP
       ��@     4�@     ��@     0�@             �@     ��@     ��@     ��@      =@     \�@      &@     `�@      &@     `p@       @     `p@       @     �C@      �?      6@              1@      �?      @      �?      @                      �?      (@             �k@      �?     �b@      �?     �`@              .@      �?       @              @      �?      @      �?      @             �R@                      @     `p@      @     �m@              7@      @      7@      �?      (@              &@      �?      @      �?      @                       @     X�@             �R@      2@      @      @      @      @      @       @      @      �?              �?              �?              �?     @Q@      ,@      ?@              C@      ,@      C@      *@      4@      @      4@       @      $@              $@       @      @       @      @                      �?      2@      $@      2@      @       @              $@      @      "@      @      @       @      @       @      �?                      @              �?             ��@     С@     �@     С@     0r@      H@      Y@      6@              :@      Y@             �S@      :@      6@      "@      6@              ,@      "@       @      @      @               @      @       @      @      @              �?      @      @      1@             p�@     �g@     h�@     @R@      C@      <@              <@      C@             И@     �F@     x�@     �F@     8�@              D@     �F@             �F@      D@             (�@             ��@     �]@     �q@     �]@     �`@     @U@      0@      6@              ,@      0@       @      $@      @      @              @      @               @      @       @      @      @       @      @       @                      @      @      �?     �]@     �O@     �X@      ,@              �?     �X@      *@      8@      @      8@                      @     �R@      @      B@      @      6@              ,@      @      ,@                      @     �C@      �?     �C@                      �?      3@     �H@      @              (@     �H@              .@      (@      A@      (@      <@      @      6@      @                      6@      "@      @      "@                      @              @      c@     �@@     �V@     �@@      0@             �R@     �@@      $@      ,@      $@                      ,@     @P@      3@      @             �M@      3@     �A@              8@      3@      @      ,@      @              �?      ,@              ,@      �?              1@      @      $@              @      @              @      @              O@             �s@                     �k@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�BX)         &                    @؆d#~��?�           c�@                           @xZ{O��?�           ܤ@                           �?��U����?�           �@������������������������       �        b           ��@                           @�b�]�?�           ��@       	                     �?������?            |@                           �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@
                           @
@�lFf�?           `{@������������������������       �        �            �n@                           �?�X-:oȤ?o             h@                           �?������?             1@������������������������       �                     *@������������������������       �                     @������������������������       �        h             f@                           @�MI8d�?�            �k@������������������������       �        t             g@                           �?�}�+r��?             C@                           �?8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     9@                           @6�i�w�?�           `�@                           @���;�f�?%           @|@                           �?Oi�8��?�            �n@������������������������       �        �            �h@������������������������       �                      G@������������������������       �        �            �i@       %                     @ �q�q�?l             e@                            �?���Hx�?3             R@������������������������       �                    �C@!       "                    �?�'�`d�?            �@@������������������������       �                      @#       $                    @ �o_��?             9@������������������������       �                     2@������������������������       �                     @������������������������       �        9             X@'       f                    �?�l��_.�?f	           �@(       Q                     @�t�"��?V           @�@)       <                    @�5;��?�            �@*       ;                    �?��T��g�?^           x�@+       :                    !@R�}e�.�?�            �q@,       /                    @ 4�"=[�?�            �n@-       .                    @����S��?I             ]@������������������������       �                     A@������������������������       �        2            �T@0       1                    !@0�ޤ��?R            @`@������������������������       �        E            @[@2       5                     �?؇���X�?             5@3       4                    @���Q��?             @������������������������       �                      @������������������������       �                     @6       7                     @      �?
             0@������������������������       �                     @8       9                    @$�q-�?             *@������������������������       �؇���X�?             @������������������������       �                     @������������������������       �                     D@������������������������       �        �            q@=       @                     @4ڗ��?\            �b@>       ?                    @��(\���?1             T@������������������������       �        .            �R@������������������������       �                     @A       P                    %@ꮃG��?+            @Q@B       O                    !@�^���U�?#            �L@C       D                    #@�z�G��?             I@������������������������       �                     @E       N                    @(���@��?            �G@F       G                    @�n_Y�K�?            �C@������������������������       �                     (@H       I                    @�����H�?             ;@������������������������       �                     @J       M                     @؇���X�?             5@K       L                     �?z�G�z�?	             .@������������������������       �      �?             @������������������������       �"pc�
�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     (@R       S                    @@܍���?�           `�@������������������������       �        �            �q@T       U                    #@�����?�             w@������������������������       �        �            �s@V       e                    !@$�q-�?#             J@W       `                    @�IєX�?"            �I@X       Y                    @P�Lt�<�?             C@������������������������       �        
             .@Z       _                    %@�nkK�?             7@[       ^                    �?@4և���?
             ,@\       ]                    @�����H�?             "@������������������������       �      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     "@a       d                    @8�Z$���?	             *@b       c                    @�<ݚ�?             "@������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @������������������������       �                     �?g       x                    �?��Ҕ��?           J�@h       q                    @L�w�=�?+            �Q@i       j                    @���c�H�?             �H@������������������������       �                    �A@k       p                     @d}h���?
             ,@l       m                    "@      �?             @������������������������       �                     �?n       o                     �?���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                      @r       s                    "@և���X�?             5@������������������������       �                      @t       w                     @p�ݯ��?
             3@u       v                     �?�z�G��?             $@������������������������       �                     @������������������������       �և���X�?             @������������������������       �                     "@y       z                    �?����I��?�           ��@������������������������       �        �           �@{       �                    @���#���?           ��@|       �                     �?�(�&��?-           �}@}       ~                    �?����1�?-            @R@������������������������       �                     @       �                    @ >�֕�?,            �Q@������������������������       �        )            �P@������������������������       �                     @�       �                    @�mX|���?            0y@�       �                    @�Ϫ�U�?�            �r@�       �                    @��+7��?.            @Q@������������������������       �        #            �I@������������������������       �                     2@�       �                    @�b(��[�?�            �l@������������������������       �        -            �T@�       �                     @�T�j��?^            @b@�       �                    �?�w��#��?%             I@������������������������       �                     �?�       �                    "@���Q �?$            �H@�       �                    @      �?             0@�       �                    !@8�Z$���?
             *@�       �                    �?�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                     @�       �                    @�eP*L��?            �@@������������������������       �                     @�       �                    �?�q�q�?             ;@������������������������       �                     @�       �                    @"pc�
�?             6@������������������������       �                     ,@�       �                    @      �?              @������������������������       �                     �?�       �                    @և���X�?             @������������������������       ����Q��?             @������������������������       �                      @�       �                    !@�q�q��?9             X@�       �                    @�Y�R_�?)            �Q@�       �                    �?�Gi����?            �B@������������������������       �        	             .@������������������������       �                     6@������������������������       �                     A@������������������������       �                     9@������������������������       �        G            @Z@�       �                    @4��A��?�           ��@�       �                     �?�	j*D�?3            �S@������������������������       �                     >@�       �                    @      �?              H@������������������������       �                     *@�       �                    @">�֕�?            �A@������������������������       �                     8@������������������������       �                     &@�       �                    @���d��?�           L�@�       �                    @��}���?�           �@������������������������       �        �            �p@�       �                    @P
�6$��?�           ��@�       �                    @���=��?�           p�@������������������������       �        �           ؆@�       �                     �?�d�����?             3@������������������������       �                     @�       �                     @      �?	             0@�       �                    "@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �        9             T@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B�       ��@     �@     �{@     j�@     @m@     `�@             ��@     @m@     @{@     �h@     @o@      "@      �?              �?      "@             �g@      o@             �n@     �g@      @      *@      @      *@                      @      f@              B@     @g@              g@      B@       @      &@       @      &@                       @      9@             �i@     �y@      G@     `y@      G@     �h@             �h@      G@                     �i@      d@      @     @P@      @     �C@              :@      @       @              2@      @      2@                      @      X@             >�@     ��@     ȋ@     p}@     X�@      g@      ~@     @S@      j@     @S@      j@     �B@     �T@      A@              A@     �T@             �_@      @     @[@              2@      @      @       @               @      @              .@      �?      @              (@      �?      @      �?      @                      D@     q@             �D@      [@      @     �R@             �R@      @             �A@      A@     �A@      6@     �A@      .@      @              @@      .@      8@      .@              (@      8@      @      @              2@      @      (@      @      @      �?      "@       @      @               @                      @              (@     �v@     �q@             �q@     �v@      @     �s@              H@      @      H@      @     �B@      �?      .@              6@      �?      *@      �?       @      �?      �?      �?      @              @              "@              &@       @      @       @      �?              @       @      @                      �?     L�@     �w@      7@     �G@      &@      C@             �A@      &@      @      @      @              �?      @       @              �?      @      �?       @              (@      "@               @      (@      @      @      @              @      @      @      "@             �@      u@     �@             ��@      u@      p@     @k@     �P@      @              @     �P@      @     �P@                      @      h@     `j@      h@     �Z@      2@     �I@             �I@      2@             �e@     �K@     �T@             �V@     �K@      1@     �@@              �?      1@      @@       @      ,@       @      &@      �?      &@      �?                      &@      �?                      @      .@      2@      @              "@      2@      @              @      2@              ,@      @      @      �?              @      @      @       @               @     �R@      6@     �H@      6@      .@      6@      .@                      6@      A@              9@                     @Z@     ��@     �]@      K@      8@      >@              8@      8@              *@      8@      &@      8@                      &@     ��@     �W@     ��@      ,@     �p@             H�@      ,@     H�@      @     ؆@              ,@      @              @      ,@       @      @       @               @      @               @                      "@              T@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK˅�hi�Bh,         @                    @|����?           c�@       -                    �?ȫ���"�?�           ��@                           �? o�ŏ�?�           ��@������������������������       �        r           ؕ@       ,                    !@:�{��x�?�           P�@                            �?�
^��S�?�           �@������������������������       �                     7@       '                    @�jF��?�           0�@	                            @      �?"            |@
                           @�R VK5�?q            @f@                           @��S�ۿ?'             N@                           @0�)AU��?$            �L@������������������������       �        #             L@������������������������       �                     �?������������������������       �                     @                           @$��9��?J            �]@                           �?,���y4�?+             S@                           @d��0u��?!             N@������������������������       �                    �G@������������������������       �                     *@������������������������       �        
             0@������������������������       �                     E@       $                    @N�?�0��?�             q@                           �?��T���?d            @b@                           @$f����?P            @]@                           @P̏����?&            �L@������������������������       �                    �E@������������������������       �        	             ,@                           @��0u���?*             N@������������������������       �                    �E@������������������������       �                     1@        #                    @V�a�� �?             =@!       "                    @ҳ�wY;�?             1@������������������������       �                     @������������������������       �                     &@������������������������       �        	             (@%       &                    @���N8�?M            �_@������������������������       �                     >@������������������������       �        =             X@(       )                    @ؗp�'ʸ?�            �h@������������������������       �        ;            �V@*       +                    @�����?F            @Z@������������������������       �        A            �W@������������������������       �                     $@������������������������       �        �            �t@.       =                     @j����b�?�            �n@/       <                    @��
ц��?M            @]@0       7                    �?p`q�q��?5            �S@1       4                    @�	j*D�?             *@2       3                    �?      �?             @������������������������       �                      @������������������������       �                      @5       6                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @8       9                    @��IF�E�?.            �P@������������������������       �                    �B@:       ;                    �?>���Rp�?             =@������������������������       �                     6@������������������������       �                     @������������������������       �                     C@>       ?                    @@w��_m�?P            �_@������������������������       �        ;             Y@������������������������       �                     ;@A       P                    @pHR�4�?|	           �@B       I                    @̠�[�?           ,�@C       H                    �?`�E���?�            @x@D       E                     @Х-��ٹ?Y            �b@������������������������       �        .            @R@F       G                    @�s�c���?+            @S@������������������������       �                      @������������������������       �        %            @Q@������������������������       �        �            �m@J       O                    @B��,-H�?           8�@K       N                    �?8��l6�?�           ؆@L       M                    @��X��?�             u@������������������������       �                     ;@������������������������       �        �            Ps@������������������������       �        �            �x@������������������������       �        G             [@Q       �                    �?Ј�^�i�?z           ��@R       _                     �?X*,�&��?S            �@S       T                    !@h�����?6             U@������������������������       �                     ;@U       ^                    !@�}�+r��?$            �L@V       ]                    %@ �Jj�G�?"            �K@W       \                    �? ���J��?            �C@X       [                    @�IєX�?             1@Y       Z                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     6@������������������������       �        	             0@������������������������       �                      @`       �                    !@8�l���?           ��@a       ~                     @�va%n�?�           ؄@b       c                    @^H���+�?�            �t@������������������������       �        B            �Z@d       }                     @�D�n���?�            `l@e       t                    @P���Q�?�            �k@f       g                    @��?^�k�?o            �e@������������������������       �        &            @P@h       s                    @���7�?I            �[@i       j                    !@�[|x��?)            �O@������������������������       �                     =@k       p                     @��hJ,�?             A@l       o                    %@R���Q�?
             4@m       n                    �?      �?              @������������������������       �և���X�?             @������������������������       �                     �?������������������������       �                     (@q       r                    %@؇���X�?             ,@������������������������       �      �?             @������������������������       �                     $@������������������������       �                     �G@u       |                    @�r����?            �F@v       y                     @��+7��?             7@w       x                    @�q�q�?             (@������������������������       �                     @������������������������       �      �?              @z       {                    @"pc�
�?             &@������������������������       �                     @������������������������       ����Q��?             @������������������������       �                     6@������������������������       �                     @       �                    @"�!���?�            �t@�       �                    �?�1��n�?w            �e@�       �                    @X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �                    @&�bi��?q            �d@������������������������       �        M            �Z@������������������������       �        $            �L@�       �                    @&� �N�?b             d@�       �                    @���c���?#             J@�       �                    !@`Ӹ����?             �F@������������������������       �                     ?@�       �                    �?؇���X�?             ,@������������������������       �      �?              @������������������������       �                     @�       �                    @����X�?             @������������������������       �                     @������������������������       �                      @�       �                    @�A�|O��??            @[@������������������������       �                     @@�       �                    @����X�?.            @S@������������������������       �                     6@������������������������       �        "            �K@������������������������       �        u            �f@�       �                    �?V�6V>�?'           ��@������������������������       �        O           ��@�       �                    @LCI�&�?�            �@�       �                     �?�g�?�           ��@�       �                    @�P�*�?+             O@������������������������       �                     B@������������������������       �                     :@�       �                    @Tb.��?i           @�@�       �                    �?L5����?�            @o@������������������������       �        =            @Y@������������������������       �        a            �b@�       �                    �?��d>�H�?�           p�@������������������������       �                     @�       �                    @ ��-�?�           P�@�       �                    �?���W���?8            �U@�       �                     @�	j*D�?	             *@�       �                    "@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                     @���;QU�?/            @R@�       �                    @���B���?             :@������������������������       �                     $@�       �                    !@     ��?             0@�       �                    @�n_Y�K�?
             *@�       �                    "@և���X�?             @������������������������       �                      @������������������������       �z�G�z�?             @�       �                    @�q�q�?             @������������������������       �                      @�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                    �G@�       �                     @����r�?�           ��@�       �                    @�#��g1�?�            �s@������������������������       �                     5@�       �                    #@� yt5��?�            Pr@�       �                    @�����?g            �e@������������������������       �        1            �U@�       �                    !@��f�{��?6            �U@������������������������       �                     �?������������������������       �        5            @U@�       �                    @ �q�q�?N             ^@�       �                    �?���<_�?L            �]@������������������������       ����Q��?             @�       �                    @�H�I���?H            @\@������������������������       �        B            �Y@������������������������       ��C��2(�?             &@������������������������       �                      @������������������������       �        �            �u@������������������������       �        D            �X@�t�bh�h,h/K ��h1��R�(KK�KK��hJ�B�       P�@     v�@     Pz@     ^�@      p@     ��@             ؕ@      p@     @�@      p@     �y@      7@             `m@     �y@      l@      l@     �R@     �Y@      @      L@      �?      L@              L@      �?              @             �Q@     �G@      =@     �G@      *@     �G@             �G@      *@              0@              E@             �b@     �^@      K@      W@      ?@     �U@      ,@     �E@             �E@      ,@              1@     �E@             �E@      1@              7@      @      &@      @              @      &@              (@              X@      >@              >@      X@              $@     @g@             �V@      $@     �W@             �W@      $@                     �t@     `d@     @T@     �O@      K@     �O@      0@      @      "@       @       @       @                       @       @      @       @                      @     �M@      @     �B@              6@      @      6@                      @              C@      Y@      ;@      Y@                      ;@     �@     `�@     �@     �a@     �w@       @     �a@       @     @R@             @Q@       @               @     @Q@             �m@              �@     �`@      �@      ;@     Ps@      ;@              ;@     Ps@             �x@                      [@     �@     �@     �|@     �}@     @T@      @      ;@              K@      @      K@      �?      C@      �?      0@      �?      @      �?      @                      �?      &@              6@              0@                       @     �w@     `}@     �w@     r@      k@     @]@             �Z@      k@      &@      j@      &@     @e@      @     @P@             @Z@      @      M@      @      =@              =@      @      1@      @      @      @      @      @      �?              (@              (@       @       @       @      $@             �G@             �C@      @      1@      @       @      @      @              @      @      "@       @      @              @       @      6@              @             @d@     �e@      O@     �[@      @      @              @      @             �L@     �Z@             �Z@     �L@              Y@     �N@     �F@      @     �E@       @      ?@              (@       @      @       @      @               @      @              @       @             �K@      K@              @@     �K@      6@              6@     �K@                     �f@     �@     @r@     ��@              �@     @r@      �@     @h@      B@      :@      B@                      :@      �@      e@     @Y@     �b@     @Y@                     �b@     ؆@      3@              @     ؆@      .@     @S@      "@      "@      @      @      @              @      @              @              Q@      @      5@      @      $@              &@      @       @      @      @      @               @      @      �?      @       @       @               @       @       @                       @      @             �G@             p�@      @     @s@      @      5@             �q@      @     �e@      �?     �U@             @U@      �?              �?     @U@             �\@      @     �\@      @      @       @      \@      �?     �Y@              $@      �?               @     �u@                     �X@�t�bubhhubehhub.